module top (
    output wire [7:0] led
);
    assign led = 8'b10101010;
endmodule
