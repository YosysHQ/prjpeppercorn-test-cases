module neorv32_cpu_cp_muldiv_9159cb8bcee7fcb95582f140960cdae72788d326
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_lsu_req,
   input  ctrl_i_lsu_rw,
   input  ctrl_i_lsu_mo_we,
   input  ctrl_i_lsu_fence,
   input  ctrl_i_lsu_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  start_i,
   input  [31:0] rs1_i,
   input  [31:0] rs2_i,
   output [31:0] res_o,
   output valid_o);
  wire [66:0] n10117_o;
  wire [41:0] ctrl;
  wire [162:0] div;
  wire [230:0] mul;
  wire n10121_o;
  wire [1:0] n10129_o;
  wire [1:0] n10132_o;
  wire n10134_o;
  wire n10135_o;
  wire n10136_o;
  wire n10137_o;
  wire n10144_o;
  wire n10146_o;
  wire n10148_o;
  wire n10149_o;
  wire n10150_o;
  wire n10151_o;
  wire n10152_o;
  wire n10153_o;
  wire n10154_o;
  wire n10155_o;
  wire n10156_o;
  wire n10157_o;
  wire n10158_o;
  wire n10159_o;
  wire n10160_o;
  wire n10161_o;
  wire n10162_o;
  wire n10163_o;
  wire n10164_o;
  wire n10165_o;
  wire n10166_o;
  wire n10167_o;
  wire n10168_o;
  wire n10169_o;
  wire n10170_o;
  wire n10171_o;
  wire n10172_o;
  wire n10173_o;
  wire n10174_o;
  wire n10175_o;
  wire n10176_o;
  wire n10177_o;
  wire n10178_o;
  wire n10179_o;
  wire n10180_o;
  wire n10181_o;
  wire n10182_o;
  wire n10183_o;
  wire n10184_o;
  wire n10185_o;
  wire n10186_o;
  wire n10187_o;
  wire n10188_o;
  wire n10189_o;
  wire n10190_o;
  wire n10191_o;
  wire n10192_o;
  wire n10193_o;
  wire n10194_o;
  wire n10195_o;
  wire n10196_o;
  wire n10197_o;
  wire n10198_o;
  wire n10199_o;
  wire n10200_o;
  wire n10201_o;
  wire n10202_o;
  wire n10203_o;
  wire n10204_o;
  wire n10205_o;
  wire n10206_o;
  wire n10207_o;
  wire n10208_o;
  wire n10209_o;
  wire n10210_o;
  wire [1:0] n10211_o;
  wire n10213_o;
  wire n10214_o;
  wire n10216_o;
  wire n10217_o;
  wire n10218_o;
  wire n10219_o;
  wire n10220_o;
  wire [31:0] n10222_o;
  wire [31:0] n10223_o;
  wire n10224_o;
  wire n10225_o;
  wire n10227_o;
  wire [1:0] n10230_o;
  wire [1:0] n10231_o;
  wire [1:0] n10232_o;
  wire [31:0] n10233_o;
  wire [31:0] n10234_o;
  wire n10235_o;
  wire n10236_o;
  wire n10238_o;
  wire [4:0] n10239_o;
  wire [4:0] n10241_o;
  wire n10249_o;
  wire n10251_o;
  wire n10253_o;
  wire n10254_o;
  wire n10255_o;
  wire n10256_o;
  wire n10257_o;
  wire n10258_o;
  wire n10259_o;
  wire n10260_o;
  wire n10261_o;
  wire n10262_o;
  wire n10263_o;
  wire [1:0] n10265_o;
  wire [1:0] n10266_o;
  wire n10268_o;
  wire n10272_o;
  wire [2:0] n10274_o;
  reg [1:0] n10275_o;
  wire [4:0] n10276_o;
  reg [4:0] n10277_o;
  reg n10278_o;
  wire [31:0] n10279_o;
  reg [31:0] n10280_o;
  wire n10281_o;
  reg n10282_o;
  wire [6:0] n10283_o;
  wire [32:0] n10284_o;
  wire [6:0] n10291_o;
  wire [32:0] n10292_o;
  wire [1:0] n10298_o;
  wire n10300_o;
  wire n10301_o;
  wire [2:0] n10304_o;
  wire n10306_o;
  wire [2:0] n10307_o;
  wire n10309_o;
  wire n10310_o;
  wire [2:0] n10311_o;
  wire n10313_o;
  wire n10314_o;
  wire [2:0] n10315_o;
  wire n10317_o;
  wire n10318_o;
  wire n10319_o;
  wire [2:0] n10322_o;
  wire n10324_o;
  wire [2:0] n10325_o;
  wire n10327_o;
  wire n10328_o;
  wire [2:0] n10329_o;
  wire n10331_o;
  wire n10332_o;
  wire n10333_o;
  wire n10336_o;
  wire n10337_o;
  wire n10338_o;
  wire n10339_o;
  wire n10342_o;
  wire n10343_o;
  wire n10344_o;
  wire n10347_o;
  wire n10352_o;
  wire n10353_o;
  wire n10354_o;
  wire n10355_o;
  wire [32:0] n10356_o;
  wire n10357_o;
  wire n10358_o;
  wire n10359_o;
  wire [32:0] n10360_o;
  wire [65:0] n10361_o;
  wire [63:0] n10364_o;
  wire [65:0] n10369_o;
  wire [32:0] n10373_o;
  wire [32:0] n10374_o;
  wire [65:0] n10375_o;
  wire [65:0] n10376_o;
  wire [65:0] n10377_o;
  wire n10381_o;
  wire n10385_o;
  wire n10386_o;
  wire n10387_o;
  wire n10388_o;
  wire [31:0] n10390_o;
  wire [31:0] n10391_o;
  wire [1:0] n10393_o;
  wire n10395_o;
  wire [1:0] n10396_o;
  wire n10398_o;
  wire n10399_o;
  wire [30:0] n10400_o;
  wire n10401_o;
  wire n10402_o;
  wire [31:0] n10403_o;
  wire n10404_o;
  wire n10405_o;
  wire [31:0] n10406_o;
  wire [30:0] n10407_o;
  wire n10408_o;
  wire [31:0] n10409_o;
  wire [31:0] n10410_o;
  wire [63:0] n10411_o;
  wire [63:0] n10412_o;
  wire [63:0] n10413_o;
  wire [63:0] n10414_o;
  wire [63:0] n10415_o;
  wire [63:0] n10418_o;
  wire [30:0] n10421_o;
  wire [31:0] n10423_o;
  wire n10424_o;
  wire [32:0] n10425_o;
  wire [31:0] n10426_o;
  wire [32:0] n10428_o;
  wire [32:0] n10429_o;
  wire [31:0] n10430_o;
  wire [2:0] n10431_o;
  wire n10433_o;
  wire [2:0] n10434_o;
  wire n10436_o;
  wire n10437_o;
  wire [31:0] n10438_o;
  wire [31:0] n10439_o;
  wire [31:0] n10440_o;
  wire [31:0] n10442_o;
  wire n10443_o;
  wire [31:0] n10444_o;
  wire [31:0] n10445_o;
  wire n10447_o;
  wire [2:0] n10448_o;
  wire [31:0] n10449_o;
  wire n10451_o;
  wire [31:0] n10452_o;
  wire n10454_o;
  wire n10456_o;
  wire n10457_o;
  wire n10459_o;
  wire n10460_o;
  wire [31:0] n10461_o;
  wire [1:0] n10462_o;
  reg [31:0] n10463_o;
  wire [31:0] n10465_o;
  reg [32:0] n10468_q;
  reg [6:0] n10469_q;
  wire [41:0] n10470_o;
  reg [63:0] n10471_q;
  reg n10472_q;
  wire [162:0] n10473_o;
  wire [65:0] n10474_o;
  wire [65:0] n10475_o;
  reg [65:0] n10476_q;
  reg [63:0] n10477_q;
  wire [230:0] n10478_o;
  assign res_o = n10465_o; //(module output)
  assign valid_o = n10301_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:58:5  */
  assign n10117_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_lsu_priv, ctrl_i_lsu_fence, ctrl_i_lsu_mo_we, ctrl_i_lsu_rw, ctrl_i_lsu_req, ctrl_i_alu_cp_trig, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:87:10  */
  assign ctrl = n10470_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:99:10  */
  assign div = n10473_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:111:10  */
  assign mul = n10478_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:119:16  */
  assign n10121_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:130:17  */
  assign n10129_o = ctrl[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:137:35  */
  assign n10132_o = n10117_o[42:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:137:48  */
  assign n10134_o = n10132_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:138:39  */
  assign n10135_o = rs1_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:138:61  */
  assign n10136_o = rs2_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:138:52  */
  assign n10137_o = n10135_o ^ n10136_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10144_o = rs2_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10146_o = 1'b0 | n10144_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10148_o = rs2_i[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10149_o = n10146_o | n10148_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10150_o = rs2_i[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10151_o = n10149_o | n10150_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10152_o = rs2_i[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10153_o = n10151_o | n10152_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10154_o = rs2_i[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10155_o = n10153_o | n10154_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10156_o = rs2_i[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10157_o = n10155_o | n10156_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10158_o = rs2_i[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10159_o = n10157_o | n10158_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10160_o = rs2_i[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10161_o = n10159_o | n10160_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10162_o = rs2_i[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10163_o = n10161_o | n10162_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10164_o = rs2_i[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10165_o = n10163_o | n10164_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10166_o = rs2_i[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10167_o = n10165_o | n10166_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10168_o = rs2_i[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10169_o = n10167_o | n10168_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10170_o = rs2_i[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10171_o = n10169_o | n10170_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10172_o = rs2_i[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10173_o = n10171_o | n10172_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10174_o = rs2_i[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10175_o = n10173_o | n10174_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10176_o = rs2_i[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10177_o = n10175_o | n10176_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10178_o = rs2_i[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10179_o = n10177_o | n10178_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10180_o = rs2_i[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10181_o = n10179_o | n10180_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10182_o = rs2_i[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10183_o = n10181_o | n10182_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10184_o = rs2_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10185_o = n10183_o | n10184_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10186_o = rs2_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10187_o = n10185_o | n10186_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10188_o = rs2_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10189_o = n10187_o | n10188_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10190_o = rs2_i[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10191_o = n10189_o | n10190_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10192_o = rs2_i[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10193_o = n10191_o | n10192_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10194_o = rs2_i[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10195_o = n10193_o | n10194_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10196_o = rs2_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10197_o = n10195_o | n10196_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10198_o = rs2_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10199_o = n10197_o | n10198_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10200_o = rs2_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10201_o = n10199_o | n10200_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10202_o = rs2_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10203_o = n10201_o | n10202_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10204_o = rs2_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10205_o = n10203_o | n10204_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10206_o = rs2_i[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10207_o = n10205_o | n10206_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10208_o = rs2_i[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10209_o = n10207_o | n10208_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:138:75  */
  assign n10210_o = n10137_o & n10209_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:139:38  */
  assign n10211_o = n10117_o[42:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:139:51  */
  assign n10213_o = n10211_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:140:38  */
  assign n10214_o = rs1_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:139:15  */
  assign n10216_o = n10213_o ? n10214_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:137:15  */
  assign n10217_o = n10134_o ? n10210_o : n10216_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:145:25  */
  assign n10218_o = rs2_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:145:47  */
  assign n10219_o = ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:145:38  */
  assign n10220_o = n10218_o & n10219_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:146:53  */
  assign n10222_o = 32'b00000000000000000000000000000000 - rs2_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:145:15  */
  assign n10223_o = n10220_o ? n10222_o : rs2_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:152:33  */
  assign n10224_o = n10117_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:152:37  */
  assign n10225_o = ~n10224_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:152:44  */
  assign n10227_o = 1'b1 & n10225_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:152:13  */
  assign n10230_o = n10227_o ? 2'b10 : 2'b01;
  assign n10231_o = ctrl[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:134:11  */
  assign n10232_o = start_i ? n10230_o : n10231_o;
  assign n10233_o = ctrl[41:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:134:11  */
  assign n10234_o = start_i ? n10223_o : n10233_o;
  assign n10235_o = div[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:134:11  */
  assign n10236_o = start_i ? n10217_o : n10235_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:132:9  */
  assign n10238_o = n10129_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:160:55  */
  assign n10239_o = ctrl[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:160:60  */
  assign n10241_o = n10239_o - 5'b00001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10249_o = ctrl[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10251_o = 1'b0 | n10249_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10253_o = ctrl[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10254_o = n10251_o | n10253_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10255_o = ctrl[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10256_o = n10254_o | n10255_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10257_o = ctrl[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10258_o = n10256_o | n10257_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n10259_o = ctrl[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n10260_o = n10258_o | n10259_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:161:37  */
  assign n10261_o = ~n10260_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:161:55  */
  assign n10262_o = n10117_o[65]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:161:44  */
  assign n10263_o = n10261_o | n10262_o;
  assign n10265_o = ctrl[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:161:11  */
  assign n10266_o = n10263_o ? 2'b10 : n10265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:159:9  */
  assign n10268_o = n10129_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:165:9  */
  assign n10272_o = n10129_o == 2'b10;
  assign n10274_o = {n10272_o, n10268_o, n10238_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:130:7  */
  always @*
    case (n10274_o)
      3'b100: n10275_o = 2'b00;
      3'b010: n10275_o = n10266_o;
      3'b001: n10275_o = n10232_o;
      default: n10275_o = 2'b00;
    endcase
  assign n10276_o = ctrl[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:130:7  */
  always @*
    case (n10274_o)
      3'b100: n10277_o = n10276_o;
      3'b010: n10277_o = n10241_o;
      3'b001: n10277_o = 5'b11110;
      default: n10277_o = n10276_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:130:7  */
  always @*
    case (n10274_o)
      3'b100: n10278_o = 1'b1;
      3'b010: n10278_o = 1'b0;
      3'b001: n10278_o = 1'b0;
      default: n10278_o = 1'b0;
    endcase
  assign n10279_o = ctrl[41:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:130:7  */
  always @*
    case (n10274_o)
      3'b100: n10280_o = n10279_o;
      3'b010: n10280_o = n10279_o;
      3'b001: n10280_o = n10234_o;
      default: n10280_o = n10279_o;
    endcase
  assign n10281_o = div[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:130:7  */
  always @*
    case (n10274_o)
      3'b100: n10282_o = n10281_o;
      3'b010: n10282_o = n10281_o;
      3'b001: n10282_o = n10236_o;
      default: n10282_o = n10281_o;
    endcase
  assign n10283_o = {n10277_o, n10275_o};
  assign n10284_o = {n10280_o, n10278_o};
  assign n10291_o = {5'b00000, 2'b00};
  assign n10292_o = {32'b00000000000000000000000000000000, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:177:29  */
  assign n10298_o = ctrl[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:177:35  */
  assign n10300_o = n10298_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:177:18  */
  assign n10301_o = n10300_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:180:42  */
  assign n10304_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:180:52  */
  assign n10306_o = n10304_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:180:76  */
  assign n10307_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:180:86  */
  assign n10309_o = n10307_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:180:65  */
  assign n10310_o = n10306_o | n10309_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:181:42  */
  assign n10311_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:181:52  */
  assign n10313_o = n10311_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:180:101  */
  assign n10314_o = n10310_o | n10313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:181:76  */
  assign n10315_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:181:86  */
  assign n10317_o = n10315_o == 3'b110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:181:65  */
  assign n10318_o = n10314_o | n10317_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:180:29  */
  assign n10319_o = n10318_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:182:42  */
  assign n10322_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:182:52  */
  assign n10324_o = n10322_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:183:42  */
  assign n10325_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:183:52  */
  assign n10327_o = n10325_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:182:65  */
  assign n10328_o = n10324_o | n10327_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:183:76  */
  assign n10329_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:183:86  */
  assign n10331_o = n10329_o == 3'b110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:183:65  */
  assign n10332_o = n10328_o | n10331_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:182:29  */
  assign n10333_o = n10332_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:186:62  */
  assign n10336_o = n10117_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:186:66  */
  assign n10337_o = ~n10336_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:186:41  */
  assign n10338_o = n10337_o & start_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:186:20  */
  assign n10339_o = n10338_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:187:62  */
  assign n10342_o = n10117_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:187:41  */
  assign n10343_o = n10342_o & start_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:187:20  */
  assign n10344_o = n10343_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:198:18  */
  assign n10347_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:203:17  */
  assign n10352_o = mul[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:204:37  */
  assign n10353_o = rs1_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:204:59  */
  assign n10354_o = ctrl[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:204:50  */
  assign n10355_o = n10353_o & n10354_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:204:74  */
  assign n10356_o = {n10355_o, rs1_i};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:205:37  */
  assign n10357_o = rs2_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:205:59  */
  assign n10358_o = ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:205:50  */
  assign n10359_o = n10357_o & n10358_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:205:74  */
  assign n10360_o = {n10359_o, rs2_i};
  assign n10361_o = {n10360_o, n10356_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:207:48  */
  assign n10364_o = mul[228:165]; // extract
  assign n10369_o = {33'b000000000000000000000000000000000, 33'b000000000000000000000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:212:22  */
  assign n10373_o = mul[131:99]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:212:34  */
  assign n10374_o = mul[164:132]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:212:28  */
  assign n10375_o = {{33{n10373_o[32]}}, n10373_o}; // sext
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:212:28  */
  assign n10376_o = {{33{n10374_o[32]}}, n10374_o}; // sext
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:212:28  */
  assign n10377_o = $signed(n10375_o) * $signed(n10376_o); // smul
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:281:18  */
  assign n10381_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:285:17  */
  assign n10385_o = div[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:286:21  */
  assign n10386_o = rs1_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:286:43  */
  assign n10387_o = ctrl[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:286:34  */
  assign n10388_o = n10386_o & n10387_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:287:49  */
  assign n10390_o = 32'b00000000000000000000000000000000 - rs1_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:286:11  */
  assign n10391_o = n10388_o ? n10390_o : rs1_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:292:21  */
  assign n10393_o = ctrl[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:292:27  */
  assign n10395_o = n10393_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:292:46  */
  assign n10396_o = ctrl[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:292:52  */
  assign n10398_o = n10396_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:292:37  */
  assign n10399_o = n10395_o | n10398_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:293:39  */
  assign n10400_o = div[64:34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:293:67  */
  assign n10401_o = div[98]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:293:56  */
  assign n10402_o = ~n10401_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:293:53  */
  assign n10403_o = {n10400_o, n10402_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:294:22  */
  assign n10404_o = div[98]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:294:27  */
  assign n10405_o = ~n10404_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:295:37  */
  assign n10406_o = div[97:66]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:297:43  */
  assign n10407_o = div[32:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:297:71  */
  assign n10408_o = div[65]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:297:57  */
  assign n10409_o = {n10407_o, n10408_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:294:11  */
  assign n10410_o = n10405_o ? n10406_o : n10409_o;
  assign n10411_o = {n10403_o, n10410_o};
  assign n10412_o = div[65:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:292:9  */
  assign n10413_o = n10399_o ? n10411_o : n10412_o;
  assign n10414_o = {n10391_o, 32'b00000000000000000000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:285:9  */
  assign n10415_o = n10385_o ? n10414_o : n10413_o;
  assign n10418_o = {32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:304:62  */
  assign n10421_o = div[32:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:304:47  */
  assign n10423_o = {1'b0, n10421_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:304:90  */
  assign n10424_o = div[65]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:304:76  */
  assign n10425_o = {n10423_o, n10424_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:304:118  */
  assign n10426_o = ctrl[41:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:304:111  */
  assign n10428_o = {1'b0, n10426_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:304:96  */
  assign n10429_o = n10425_o - n10428_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:307:22  */
  assign n10430_o = div[65:34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:307:44  */
  assign n10431_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:307:54  */
  assign n10433_o = n10431_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:307:77  */
  assign n10434_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:307:87  */
  assign n10436_o = n10434_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:307:66  */
  assign n10437_o = n10433_o | n10436_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:307:31  */
  assign n10438_o = n10437_o ? n10430_o : n10439_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:307:109  */
  assign n10439_o = div[33:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:308:53  */
  assign n10440_o = div[130:99]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:308:38  */
  assign n10442_o = 32'b00000000000000000000000000000000 - n10440_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:308:71  */
  assign n10443_o = div[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:308:61  */
  assign n10444_o = n10443_o ? n10442_o : n10445_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:308:96  */
  assign n10445_o = div[130:99]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:328:14  */
  assign n10447_o = ctrl[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:329:19  */
  assign n10448_o = n10117_o[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:331:28  */
  assign n10449_o = mul[32:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:330:9  */
  assign n10451_o = n10448_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:333:28  */
  assign n10452_o = mul[64:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:332:9  */
  assign n10454_o = n10448_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:332:24  */
  assign n10456_o = n10448_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:332:24  */
  assign n10457_o = n10454_o | n10456_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:332:38  */
  assign n10459_o = n10448_o == 3'b011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:332:38  */
  assign n10460_o = n10457_o | n10459_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:335:24  */
  assign n10461_o = div[162:131]; // extract
  assign n10462_o = {n10460_o, n10451_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:329:7  */
  always @*
    case (n10462_o)
      2'b10: n10463_o = n10452_o;
      2'b01: n10463_o = n10449_o;
      default: n10463_o = n10461_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:328:5  */
  assign n10465_o = n10447_o ? n10463_o : 32'b00000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:125:5  */
  always @(posedge clk_i or posedge n10121_o)
    if (n10121_o)
      n10468_q <= n10292_o;
    else
      n10468_q <= n10284_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:125:5  */
  always @(posedge clk_i or posedge n10121_o)
    if (n10121_o)
      n10469_q <= n10291_o;
    else
      n10469_q <= n10283_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:119:5  */
  assign n10470_o = {n10468_q, n10333_o, n10319_o, n10469_q};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:284:7  */
  always @(posedge clk_i or posedge n10381_o)
    if (n10381_o)
      n10471_q <= n10418_o;
    else
      n10471_q <= n10415_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:125:5  */
  always @(posedge clk_i or posedge n10121_o)
    if (n10121_o)
      n10472_q <= 1'b0;
    else
      n10472_q <= n10282_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:119:5  */
  assign n10473_o = {n10444_o, n10438_o, n10429_o, n10471_q, n10472_q, n10344_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:202:7  */
  assign n10474_o = mul[164:99]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:202:7  */
  assign n10475_o = n10352_o ? n10361_o : n10474_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:202:7  */
  always @(posedge clk_i or posedge n10347_o)
    if (n10347_o)
      n10476_q <= n10369_o;
    else
      n10476_q <= n10475_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:202:7  */
  always @(posedge clk_i or posedge n10347_o)
    if (n10347_o)
      n10477_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n10477_q <= n10364_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_muldiv.vhd:198:7  */
  assign n10478_o = {n10377_o, n10476_q, 1'b0, 33'b000000000000000000000000000000000, n10477_q, n10339_o};
endmodule

module neorv32_cpu_cp_shifter_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_lsu_req,
   input  ctrl_i_lsu_rw,
   input  ctrl_i_lsu_mo_we,
   input  ctrl_i_lsu_fence,
   input  ctrl_i_lsu_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  start_i,
   input  [31:0] rs1_i,
   input  [4:0] shamt_i,
   output [31:0] res_o,
   output valid_o);
  wire [66:0] n9815_o;
  wire [191:0] bs_level;
  wire bs_start;
  wire [31:0] bs_result;
  wire n9819_o;
  wire n9820_o;
  wire n9828_o;
  wire n9831_o;
  wire n9833_o;
  wire n9835_o;
  wire n9837_o;
  wire n9839_o;
  wire n9841_o;
  wire n9843_o;
  wire n9845_o;
  wire n9847_o;
  wire n9849_o;
  wire n9851_o;
  wire n9853_o;
  wire n9855_o;
  wire n9857_o;
  wire n9859_o;
  wire n9861_o;
  wire n9863_o;
  wire n9865_o;
  wire n9867_o;
  wire n9869_o;
  wire n9871_o;
  wire n9873_o;
  wire n9875_o;
  wire n9877_o;
  wire n9879_o;
  wire n9881_o;
  wire n9883_o;
  wire n9885_o;
  wire n9887_o;
  wire n9889_o;
  wire n9891_o;
  wire [31:0] n9892_o;
  wire [31:0] n9894_o;
  wire n9896_o;
  wire n9897_o;
  wire n9898_o;
  wire n9899_o;
  wire n9900_o;
  wire n9901_o;
  wire n9902_o;
  wire n9903_o;
  wire n9904_o;
  wire n9905_o;
  wire n9906_o;
  wire n9907_o;
  wire n9908_o;
  wire n9909_o;
  wire n9910_o;
  wire n9911_o;
  wire n9912_o;
  wire n9913_o;
  wire n9914_o;
  wire n9915_o;
  wire n9916_o;
  wire n9917_o;
  wire n9918_o;
  wire n9919_o;
  wire n9920_o;
  wire n9921_o;
  wire n9922_o;
  wire n9923_o;
  wire n9924_o;
  wire n9925_o;
  wire n9926_o;
  wire n9927_o;
  wire n9928_o;
  wire n9929_o;
  wire n9930_o;
  wire n9931_o;
  wire n9932_o;
  wire n9933_o;
  wire n9934_o;
  wire n9935_o;
  wire n9936_o;
  wire n9937_o;
  wire n9938_o;
  wire n9939_o;
  wire n9940_o;
  wire n9941_o;
  wire n9942_o;
  wire n9943_o;
  wire n9944_o;
  wire [3:0] n9945_o;
  wire [3:0] n9946_o;
  wire [3:0] n9947_o;
  wire [3:0] n9948_o;
  wire [15:0] n9949_o;
  wire [15:0] n9950_o;
  wire [31:0] n9951_o;
  wire [31:0] n9952_o;
  wire [31:0] n9953_o;
  wire n9954_o;
  wire n9955_o;
  wire n9956_o;
  wire n9957_o;
  wire n9958_o;
  wire n9959_o;
  wire n9960_o;
  wire n9961_o;
  wire n9962_o;
  wire n9963_o;
  wire n9964_o;
  wire n9965_o;
  wire n9966_o;
  wire n9967_o;
  wire n9968_o;
  wire n9969_o;
  wire n9970_o;
  wire n9971_o;
  wire n9972_o;
  wire n9973_o;
  wire n9974_o;
  wire n9975_o;
  wire n9976_o;
  wire n9977_o;
  wire n9978_o;
  wire [3:0] n9979_o;
  wire [3:0] n9980_o;
  wire [7:0] n9981_o;
  wire [23:0] n9982_o;
  wire [31:0] n9983_o;
  wire [31:0] n9984_o;
  wire [31:0] n9985_o;
  wire n9986_o;
  wire n9987_o;
  wire n9988_o;
  wire n9989_o;
  wire n9990_o;
  wire n9991_o;
  wire n9992_o;
  wire n9993_o;
  wire n9994_o;
  wire n9995_o;
  wire n9996_o;
  wire n9997_o;
  wire n9998_o;
  wire [3:0] n9999_o;
  wire [27:0] n10000_o;
  wire [31:0] n10001_o;
  wire [31:0] n10002_o;
  wire [31:0] n10003_o;
  wire n10004_o;
  wire n10005_o;
  wire n10006_o;
  wire n10007_o;
  wire n10008_o;
  wire n10009_o;
  wire n10010_o;
  wire [1:0] n10011_o;
  wire [29:0] n10012_o;
  wire [31:0] n10013_o;
  wire [31:0] n10014_o;
  wire [31:0] n10015_o;
  wire n10016_o;
  wire n10017_o;
  wire n10018_o;
  wire n10019_o;
  wire [30:0] n10020_o;
  wire [31:0] n10021_o;
  wire [31:0] n10022_o;
  wire [31:0] n10023_o;
  wire n10026_o;
  wire [31:0] n10028_o;
  wire n10037_o;
  wire [31:0] n10038_o;
  wire n10045_o;
  wire n10048_o;
  wire n10050_o;
  wire n10052_o;
  wire n10054_o;
  wire n10056_o;
  wire n10058_o;
  wire n10060_o;
  wire n10062_o;
  wire n10064_o;
  wire n10066_o;
  wire n10068_o;
  wire n10070_o;
  wire n10072_o;
  wire n10074_o;
  wire n10076_o;
  wire n10078_o;
  wire n10080_o;
  wire n10082_o;
  wire n10084_o;
  wire n10086_o;
  wire n10088_o;
  wire n10090_o;
  wire n10092_o;
  wire n10094_o;
  wire n10096_o;
  wire n10098_o;
  wire n10100_o;
  wire n10102_o;
  wire n10104_o;
  wire n10106_o;
  wire n10108_o;
  wire [31:0] n10109_o;
  wire n10110_o;
  wire n10111_o;
  wire [31:0] n10112_o;
  wire [191:0] n10114_o;
  reg n10115_q;
  reg [31:0] n10116_q;
  assign res_o = n10038_o; //(module output)
  assign valid_o = start_i; //(module output)
  assign n9815_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_lsu_priv, ctrl_i_lsu_fence, ctrl_i_lsu_mo_we, ctrl_i_lsu_rw, ctrl_i_lsu_req, ctrl_i_alu_cp_trig, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:77:10  */
  assign bs_level = n10114_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:78:10  */
  assign bs_start = n10115_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:79:10  */
  assign bs_result = n10116_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:135:27  */
  assign n9819_o = n9815_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:135:31  */
  assign n9820_o = ~n9819_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9828_o = rs1_i[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9831_o = rs1_i[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9833_o = rs1_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9835_o = rs1_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9837_o = rs1_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9839_o = rs1_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9841_o = rs1_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9843_o = rs1_i[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9845_o = rs1_i[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9847_o = rs1_i[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9849_o = rs1_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9851_o = rs1_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9853_o = rs1_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9855_o = rs1_i[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9857_o = rs1_i[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9859_o = rs1_i[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9861_o = rs1_i[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9863_o = rs1_i[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9865_o = rs1_i[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9867_o = rs1_i[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9869_o = rs1_i[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9871_o = rs1_i[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9873_o = rs1_i[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9875_o = rs1_i[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9877_o = rs1_i[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9879_o = rs1_i[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9881_o = rs1_i[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9883_o = rs1_i[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9885_o = rs1_i[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9887_o = rs1_i[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9889_o = rs1_i[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n9891_o = rs1_i[31]; // extract
  assign n9892_o = {n9828_o, n9831_o, n9833_o, n9835_o, n9837_o, n9839_o, n9841_o, n9843_o, n9845_o, n9847_o, n9849_o, n9851_o, n9853_o, n9855_o, n9857_o, n9859_o, n9861_o, n9863_o, n9865_o, n9867_o, n9869_o, n9871_o, n9873_o, n9875_o, n9877_o, n9879_o, n9881_o, n9883_o, n9885_o, n9887_o, n9889_o, n9891_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:135:7  */
  assign n9894_o = n9820_o ? n9892_o : rs1_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:20  */
  assign n9896_o = shamt_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9897_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9898_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9899_o = n9897_o & n9898_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9900_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9901_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9902_o = n9900_o & n9901_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9903_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9904_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9905_o = n9903_o & n9904_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9906_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9907_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9908_o = n9906_o & n9907_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9909_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9910_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9911_o = n9909_o & n9910_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9912_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9913_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9914_o = n9912_o & n9913_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9915_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9916_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9917_o = n9915_o & n9916_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9918_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9919_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9920_o = n9918_o & n9919_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9921_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9922_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9923_o = n9921_o & n9922_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9924_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9925_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9926_o = n9924_o & n9925_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9927_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9928_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9929_o = n9927_o & n9928_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9930_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9931_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9932_o = n9930_o & n9931_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9933_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9934_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9935_o = n9933_o & n9934_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9936_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9937_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9938_o = n9936_o & n9937_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9939_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9940_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9941_o = n9939_o & n9940_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9942_o = bs_level[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9943_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9944_o = n9942_o & n9943_o;
  assign n9945_o = {n9899_o, n9902_o, n9905_o, n9908_o};
  assign n9946_o = {n9911_o, n9914_o, n9917_o, n9920_o};
  assign n9947_o = {n9923_o, n9926_o, n9929_o, n9932_o};
  assign n9948_o = {n9935_o, n9938_o, n9941_o, n9944_o};
  assign n9949_o = {n9945_o, n9946_o, n9947_o, n9948_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:144:66  */
  assign n9950_o = bs_level[191:176]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:146:34  */
  assign n9951_o = bs_level[191:160]; // extract
  assign n9952_o = {n9949_o, n9950_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:9  */
  assign n9953_o = n9896_o ? n9952_o : n9951_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:20  */
  assign n9954_o = shamt_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9955_o = bs_level[159]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9956_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9957_o = n9955_o & n9956_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9958_o = bs_level[159]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9959_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9960_o = n9958_o & n9959_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9961_o = bs_level[159]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9962_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9963_o = n9961_o & n9962_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9964_o = bs_level[159]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9965_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9966_o = n9964_o & n9965_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9967_o = bs_level[159]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9968_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9969_o = n9967_o & n9968_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9970_o = bs_level[159]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9971_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9972_o = n9970_o & n9971_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9973_o = bs_level[159]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9974_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9975_o = n9973_o & n9974_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9976_o = bs_level[159]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9977_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9978_o = n9976_o & n9977_o;
  assign n9979_o = {n9957_o, n9960_o, n9963_o, n9966_o};
  assign n9980_o = {n9969_o, n9972_o, n9975_o, n9978_o};
  assign n9981_o = {n9979_o, n9980_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:144:66  */
  assign n9982_o = bs_level[159:136]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:146:34  */
  assign n9983_o = bs_level[159:128]; // extract
  assign n9984_o = {n9981_o, n9982_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:9  */
  assign n9985_o = n9954_o ? n9984_o : n9983_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:20  */
  assign n9986_o = shamt_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9987_o = bs_level[127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9988_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9989_o = n9987_o & n9988_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9990_o = bs_level[127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9991_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9992_o = n9990_o & n9991_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9993_o = bs_level[127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9994_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9995_o = n9993_o & n9994_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n9996_o = bs_level[127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n9997_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n9998_o = n9996_o & n9997_o;
  assign n9999_o = {n9989_o, n9992_o, n9995_o, n9998_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:144:66  */
  assign n10000_o = bs_level[127:100]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:146:34  */
  assign n10001_o = bs_level[127:96]; // extract
  assign n10002_o = {n9999_o, n10000_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:9  */
  assign n10003_o = n9986_o ? n10002_o : n10001_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:20  */
  assign n10004_o = shamt_i[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n10005_o = bs_level[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n10006_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n10007_o = n10005_o & n10006_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n10008_o = bs_level[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n10009_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n10010_o = n10008_o & n10009_o;
  assign n10011_o = {n10007_o, n10010_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:144:66  */
  assign n10012_o = bs_level[95:66]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:146:34  */
  assign n10013_o = bs_level[95:64]; // extract
  assign n10014_o = {n10011_o, n10012_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:9  */
  assign n10015_o = n10004_o ? n10014_o : n10013_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:20  */
  assign n10016_o = shamt_i[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:78  */
  assign n10017_o = bs_level[63]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:108  */
  assign n10018_o = n9815_o[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:143:87  */
  assign n10019_o = n10017_o & n10018_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:144:66  */
  assign n10020_o = bs_level[63:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:146:34  */
  assign n10021_o = bs_level[63:32]; // extract
  assign n10022_o = {n10019_o, n10020_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:142:9  */
  assign n10023_o = n10016_o ? n10022_o : n10021_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:154:18  */
  assign n10026_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:159:30  */
  assign n10028_o = bs_level[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:164:45  */
  assign n10037_o = ~bs_start;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:164:30  */
  assign n10038_o = n10037_o ? 32'b00000000000000000000000000000000 : n10112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10045_o = bs_result[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10048_o = bs_result[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10050_o = bs_result[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10052_o = bs_result[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10054_o = bs_result[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10056_o = bs_result[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10058_o = bs_result[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10060_o = bs_result[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10062_o = bs_result[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10064_o = bs_result[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10066_o = bs_result[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10068_o = bs_result[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10070_o = bs_result[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10072_o = bs_result[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10074_o = bs_result[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10076_o = bs_result[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10078_o = bs_result[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10080_o = bs_result[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10082_o = bs_result[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10084_o = bs_result[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10086_o = bs_result[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10088_o = bs_result[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10090_o = bs_result[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10092_o = bs_result[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10094_o = bs_result[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10096_o = bs_result[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10098_o = bs_result[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10100_o = bs_result[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10102_o = bs_result[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10104_o = bs_result[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10106_o = bs_result[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1096:42  */
  assign n10108_o = bs_result[31]; // extract
  assign n10109_o = {n10045_o, n10048_o, n10050_o, n10052_o, n10054_o, n10056_o, n10058_o, n10060_o, n10062_o, n10064_o, n10066_o, n10068_o, n10070_o, n10072_o, n10074_o, n10076_o, n10078_o, n10080_o, n10082_o, n10084_o, n10086_o, n10088_o, n10090_o, n10092_o, n10094_o, n10096_o, n10098_o, n10100_o, n10102_o, n10104_o, n10106_o, n10108_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:165:57  */
  assign n10110_o = n9815_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:165:61  */
  assign n10111_o = ~n10110_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:164:52  */
  assign n10112_o = n10111_o ? n10109_o : bs_result;
  assign n10114_o = {n9894_o, n9953_o, n9985_o, n10003_o, n10015_o, n10023_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:157:7  */
  always @(posedge clk_i or posedge n10026_o)
    if (n10026_o)
      n10115_q <= 1'b0;
    else
      n10115_q <= start_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_cp_shifter.vhd:157:7  */
  always @(posedge clk_i or posedge n10026_o)
    if (n10026_o)
      n10116_q <= 32'b00000000000000000000000000000000;
    else
      n10116_q <= n10028_o;
endmodule

module neorv32_cpu_decompressor
  (input  [15:0] ci_instr16_i,
   output [31:0] ci_instr32_o);
  wire [20:0] imm20;
  wire [12:0] imm12;
  wire illegal;
  wire [31:0] decoded;
  wire n8990_o;
  wire n8991_o;
  wire n8992_o;
  wire n8993_o;
  wire n8994_o;
  wire n8995_o;
  wire n8996_o;
  wire n8997_o;
  wire n8998_o;
  wire n8999_o;
  wire n9000_o;
  wire n9001_o;
  wire n9002_o;
  wire n9003_o;
  wire n9004_o;
  wire n9005_o;
  wire n9006_o;
  wire n9007_o;
  wire n9008_o;
  wire n9009_o;
  wire [3:0] n9010_o;
  wire [3:0] n9011_o;
  wire [1:0] n9012_o;
  wire [9:0] n9013_o;
  wire n9015_o;
  wire n9016_o;
  wire n9017_o;
  wire n9018_o;
  wire n9019_o;
  wire n9020_o;
  wire n9021_o;
  wire n9022_o;
  wire n9023_o;
  wire n9024_o;
  wire n9025_o;
  wire n9026_o;
  wire [3:0] n9027_o;
  wire [4:0] n9028_o;
  wire [1:0] n9030_o;
  wire [2:0] n9031_o;
  wire [2:0] n9034_o;
  wire [4:0] n9036_o;
  localparam [11:0] n9038_o = 12'b000000000000;
  wire n9043_o;
  wire n9045_o;
  wire n9047_o;
  wire n9049_o;
  wire n9051_o;
  wire n9053_o;
  wire n9055_o;
  wire n9057_o;
  wire [1:0] n9058_o;
  wire [7:0] n9059_o;
  wire n9061_o;
  wire n9064_o;
  wire n9066_o;
  localparam [1:0] n9068_o = 2'b00;
  wire n9069_o;
  wire n9070_o;
  wire n9071_o;
  wire n9072_o;
  wire n9073_o;
  localparam [4:0] n9074_o = 5'b00000;
  wire [2:0] n9076_o;
  wire [4:0] n9078_o;
  wire [2:0] n9079_o;
  wire [4:0] n9081_o;
  wire n9083_o;
  wire n9086_o;
  wire n9087_o;
  wire n9088_o;
  wire n9089_o;
  wire n9090_o;
  localparam [4:0] n9091_o = 5'b00000;
  wire [2:0] n9093_o;
  wire [4:0] n9095_o;
  wire [2:0] n9096_o;
  wire [4:0] n9098_o;
  wire n9100_o;
  wire [2:0] n9101_o;
  reg n9104_o;
  reg [6:0] n9106_o;
  wire [1:0] n9107_o;
  wire [1:0] n9108_o;
  reg [1:0] n9110_o;
  wire n9111_o;
  wire n9112_o;
  reg n9114_o;
  wire n9115_o;
  wire n9116_o;
  reg n9118_o;
  wire n9119_o;
  wire n9120_o;
  reg n9122_o;
  reg [2:0] n9124_o;
  reg [4:0] n9126_o;
  wire n9127_o;
  wire n9128_o;
  reg n9130_o;
  wire n9131_o;
  wire n9132_o;
  reg n9134_o;
  wire n9135_o;
  reg n9137_o;
  wire n9138_o;
  reg n9140_o;
  wire n9141_o;
  reg n9143_o;
  reg n9145_o;
  reg n9147_o;
  wire n9148_o;
  wire n9149_o;
  reg n9151_o;
  wire n9152_o;
  wire n9153_o;
  reg n9155_o;
  wire n9156_o;
  wire n9157_o;
  reg n9159_o;
  wire [1:0] n9160_o;
  wire [1:0] n9161_o;
  reg [1:0] n9163_o;
  wire n9165_o;
  wire [2:0] n9166_o;
  wire n9167_o;
  wire [4:0] n9170_o;
  wire [7:0] n9172_o;
  wire n9173_o;
  wire [9:0] n9174_o;
  wire n9175_o;
  wire n9177_o;
  wire n9179_o;
  wire n9180_o;
  wire n9181_o;
  wire n9182_o;
  wire [2:0] n9185_o;
  wire [2:0] n9187_o;
  wire [4:0] n9189_o;
  localparam [4:0] n9190_o = 5'b00000;
  wire n9191_o;
  wire [3:0] n9192_o;
  wire [5:0] n9193_o;
  wire n9194_o;
  wire n9196_o;
  wire n9198_o;
  wire n9199_o;
  wire [4:0] n9201_o;
  wire n9202_o;
  wire n9203_o;
  wire n9204_o;
  wire n9205_o;
  wire n9206_o;
  wire n9207_o;
  wire n9208_o;
  wire n9209_o;
  wire n9210_o;
  wire n9211_o;
  wire n9212_o;
  wire n9213_o;
  wire [3:0] n9214_o;
  wire [3:0] n9215_o;
  wire [3:0] n9216_o;
  wire [11:0] n9217_o;
  wire n9218_o;
  wire n9220_o;
  wire n9222_o;
  wire n9224_o;
  wire n9226_o;
  wire n9228_o;
  wire [5:0] n9229_o;
  wire n9231_o;
  wire [4:0] n9232_o;
  wire n9234_o;
  wire n9238_o;
  wire n9239_o;
  wire n9240_o;
  wire n9241_o;
  wire n9242_o;
  wire n9243_o;
  wire n9244_o;
  wire n9245_o;
  wire n9246_o;
  wire n9247_o;
  wire n9248_o;
  wire n9249_o;
  wire [3:0] n9250_o;
  wire [3:0] n9251_o;
  wire [3:0] n9252_o;
  wire [11:0] n9253_o;
  wire n9262_o;
  wire n9264_o;
  wire n9266_o;
  wire n9268_o;
  wire n9270_o;
  wire n9272_o;
  wire [1:0] n9273_o;
  wire [4:0] n9275_o;
  wire n9276_o;
  wire n9277_o;
  wire n9278_o;
  wire n9279_o;
  wire n9280_o;
  wire n9281_o;
  wire n9282_o;
  wire n9283_o;
  wire n9284_o;
  wire n9285_o;
  wire n9286_o;
  wire n9287_o;
  wire n9288_o;
  wire n9289_o;
  wire n9290_o;
  wire n9291_o;
  wire n9292_o;
  wire n9293_o;
  wire n9294_o;
  wire n9295_o;
  wire [3:0] n9296_o;
  wire [3:0] n9297_o;
  wire [3:0] n9298_o;
  wire [3:0] n9299_o;
  wire [3:0] n9300_o;
  wire [15:0] n9301_o;
  wire [19:0] n9302_o;
  wire n9303_o;
  wire n9305_o;
  wire n9307_o;
  wire n9309_o;
  wire n9311_o;
  wire n9313_o;
  wire [13:0] n9314_o;
  wire [31:0] n9315_o;
  wire [31:0] n9316_o;
  wire [31:0] n9317_o;
  wire [4:0] n9318_o;
  wire n9320_o;
  wire n9321_o;
  wire n9322_o;
  wire n9323_o;
  wire n9326_o;
  wire n9328_o;
  wire [4:0] n9329_o;
  wire [4:0] n9330_o;
  wire n9331_o;
  wire n9332_o;
  wire n9333_o;
  wire n9334_o;
  wire n9335_o;
  wire n9336_o;
  wire n9337_o;
  wire n9338_o;
  wire n9339_o;
  wire n9340_o;
  wire n9341_o;
  wire n9342_o;
  wire [3:0] n9343_o;
  wire [3:0] n9344_o;
  wire [3:0] n9345_o;
  wire [11:0] n9346_o;
  wire n9347_o;
  wire n9349_o;
  wire n9351_o;
  wire n9353_o;
  wire n9355_o;
  wire n9357_o;
  wire [5:0] n9358_o;
  wire n9360_o;
  wire [2:0] n9361_o;
  wire [4:0] n9363_o;
  wire [2:0] n9364_o;
  wire [4:0] n9366_o;
  wire [2:0] n9367_o;
  wire [4:0] n9369_o;
  wire [1:0] n9370_o;
  wire n9371_o;
  wire n9372_o;
  wire [6:0] n9375_o;
  wire n9377_o;
  wire n9378_o;
  wire n9379_o;
  wire n9380_o;
  wire n9381_o;
  wire n9382_o;
  wire n9385_o;
  wire n9387_o;
  wire n9389_o;
  wire n9390_o;
  wire n9392_o;
  wire n9393_o;
  wire n9394_o;
  wire n9395_o;
  wire n9396_o;
  wire n9397_o;
  wire n9398_o;
  wire n9399_o;
  wire n9400_o;
  wire n9401_o;
  wire n9402_o;
  wire n9403_o;
  wire [3:0] n9404_o;
  wire [3:0] n9405_o;
  wire [3:0] n9406_o;
  wire [11:0] n9407_o;
  wire n9408_o;
  wire n9410_o;
  wire n9412_o;
  wire n9414_o;
  wire n9416_o;
  wire n9418_o;
  wire [5:0] n9419_o;
  wire n9421_o;
  wire [1:0] n9423_o;
  wire n9426_o;
  wire n9430_o;
  wire n9434_o;
  wire [2:0] n9436_o;
  reg [2:0] n9437_o;
  reg [6:0] n9438_o;
  wire n9439_o;
  wire n9442_o;
  wire [1:0] n9443_o;
  reg n9445_o;
  reg [6:0] n9446_o;
  reg [2:0] n9447_o;
  wire n9448_o;
  reg n9449_o;
  wire n9450_o;
  reg n9451_o;
  wire n9452_o;
  reg n9453_o;
  wire n9454_o;
  reg n9455_o;
  wire n9456_o;
  reg n9457_o;
  wire n9458_o;
  wire n9459_o;
  reg n9460_o;
  wire [5:0] n9461_o;
  wire [5:0] n9462_o;
  reg [5:0] n9463_o;
  wire [4:0] n9468_o;
  reg n9470_o;
  wire [6:0] n9471_o;
  reg [6:0] n9472_o;
  wire n9473_o;
  wire n9474_o;
  wire n9475_o;
  wire n9476_o;
  wire n9477_o;
  reg n9478_o;
  wire [3:0] n9479_o;
  wire [3:0] n9480_o;
  wire [3:0] n9481_o;
  wire [3:0] n9482_o;
  wire [3:0] n9483_o;
  reg [3:0] n9484_o;
  wire [2:0] n9485_o;
  wire [2:0] n9486_o;
  reg [2:0] n9487_o;
  wire [4:0] n9488_o;
  wire [4:0] n9489_o;
  reg [4:0] n9490_o;
  wire n9491_o;
  wire n9492_o;
  reg n9493_o;
  wire n9494_o;
  wire n9495_o;
  wire n9496_o;
  reg n9497_o;
  wire n9498_o;
  wire n9499_o;
  wire n9500_o;
  reg n9501_o;
  wire n9502_o;
  wire n9503_o;
  wire n9504_o;
  reg n9505_o;
  wire n9506_o;
  wire n9507_o;
  wire n9508_o;
  reg n9509_o;
  wire n9510_o;
  wire n9511_o;
  wire n9512_o;
  reg n9513_o;
  wire [4:0] n9514_o;
  wire [4:0] n9515_o;
  wire [4:0] n9516_o;
  wire [4:0] n9517_o;
  wire [4:0] n9518_o;
  wire [4:0] n9519_o;
  reg [4:0] n9520_o;
  wire n9521_o;
  wire n9522_o;
  wire n9523_o;
  wire n9524_o;
  reg n9525_o;
  wire n9527_o;
  wire [2:0] n9528_o;
  wire [4:0] n9529_o;
  wire [4:0] n9530_o;
  localparam [6:0] n9532_o = 7'b0000000;
  wire n9533_o;
  wire n9534_o;
  wire n9535_o;
  wire n9536_o;
  wire n9537_o;
  wire n9538_o;
  wire n9541_o;
  wire n9543_o;
  localparam [1:0] n9544_o = 2'b00;
  wire n9545_o;
  wire n9546_o;
  wire n9547_o;
  wire n9548_o;
  wire n9549_o;
  wire n9550_o;
  wire [4:0] n9553_o;
  wire n9554_o;
  wire [4:0] n9555_o;
  wire n9557_o;
  wire n9558_o;
  wire n9561_o;
  wire n9563_o;
  wire n9565_o;
  wire n9566_o;
  wire n9568_o;
  wire n9569_o;
  wire n9570_o;
  wire n9571_o;
  wire n9572_o;
  wire n9573_o;
  wire [4:0] n9576_o;
  wire n9577_o;
  wire n9580_o;
  wire n9582_o;
  wire n9584_o;
  wire n9585_o;
  wire n9586_o;
  wire n9587_o;
  wire [4:0] n9588_o;
  wire n9590_o;
  wire [4:0] n9592_o;
  wire [4:0] n9594_o;
  wire n9596_o;
  wire [4:0] n9597_o;
  wire n9599_o;
  wire n9600_o;
  wire n9603_o;
  wire [4:0] n9605_o;
  wire [4:0] n9607_o;
  wire [4:0] n9608_o;
  wire n9610_o;
  wire n9613_o;
  wire n9614_o;
  wire [24:0] n9615_o;
  wire [11:0] n9616_o;
  wire [11:0] n9617_o;
  wire [11:0] n9618_o;
  wire [2:0] n9619_o;
  wire [2:0] n9621_o;
  wire [4:0] n9622_o;
  wire [4:0] n9623_o;
  wire [4:0] n9624_o;
  wire [4:0] n9626_o;
  wire [4:0] n9627_o;
  wire n9629_o;
  wire [4:0] n9630_o;
  wire n9632_o;
  wire [4:0] n9635_o;
  wire [11:0] n9637_o;
  wire [6:0] n9638_o;
  wire [6:0] n9639_o;
  wire [4:0] n9640_o;
  wire [4:0] n9642_o;
  wire [4:0] n9644_o;
  wire [11:0] n9646_o;
  wire [4:0] n9648_o;
  wire [4:0] n9649_o;
  wire [4:0] n9650_o;
  wire [24:0] n9651_o;
  wire [11:0] n9652_o;
  wire [16:0] n9653_o;
  wire [11:0] n9654_o;
  wire [11:0] n9655_o;
  wire [2:0] n9656_o;
  wire [2:0] n9658_o;
  wire [9:0] n9659_o;
  wire [9:0] n9660_o;
  wire [9:0] n9661_o;
  wire [6:0] n9662_o;
  wire [6:0] n9664_o;
  wire n9666_o;
  wire [31:0] n9667_o;
  wire [24:0] n9668_o;
  wire [24:0] n9669_o;
  wire [24:0] n9670_o;
  wire [6:0] n9671_o;
  wire [6:0] n9673_o;
  wire n9675_o;
  wire [3:0] n9676_o;
  reg n9678_o;
  wire [6:0] n9679_o;
  reg [6:0] n9681_o;
  wire [1:0] n9682_o;
  wire [1:0] n9683_o;
  wire [1:0] n9684_o;
  reg [1:0] n9686_o;
  wire n9687_o;
  wire n9688_o;
  wire n9689_o;
  reg n9691_o;
  wire n9692_o;
  wire n9693_o;
  wire n9694_o;
  reg n9696_o;
  wire n9697_o;
  wire n9698_o;
  wire n9699_o;
  reg n9701_o;
  wire [2:0] n9702_o;
  reg [2:0] n9704_o;
  wire [4:0] n9705_o;
  reg [4:0] n9707_o;
  wire n9708_o;
  wire n9709_o;
  wire n9710_o;
  reg n9712_o;
  wire n9713_o;
  wire n9714_o;
  wire n9715_o;
  reg n9717_o;
  wire n9718_o;
  wire n9719_o;
  reg n9721_o;
  wire n9722_o;
  wire n9723_o;
  reg n9725_o;
  wire n9726_o;
  wire n9727_o;
  reg n9729_o;
  wire n9730_o;
  wire n9731_o;
  reg n9733_o;
  wire n9734_o;
  wire n9735_o;
  reg n9737_o;
  wire n9738_o;
  wire n9739_o;
  reg n9741_o;
  wire [3:0] n9742_o;
  wire [3:0] n9743_o;
  reg [3:0] n9745_o;
  wire [1:0] n9746_o;
  reg n9747_o;
  reg [6:0] n9749_o;
  wire n9750_o;
  wire n9751_o;
  reg n9752_o;
  wire n9753_o;
  wire n9754_o;
  wire n9755_o;
  reg n9756_o;
  wire n9757_o;
  reg n9758_o;
  wire n9759_o;
  reg n9760_o;
  wire n9761_o;
  reg n9762_o;
  reg [2:0] n9763_o;
  reg [4:0] n9764_o;
  reg n9765_o;
  reg n9766_o;
  reg n9767_o;
  reg n9768_o;
  reg n9769_o;
  reg n9770_o;
  wire n9771_o;
  reg n9772_o;
  wire n9773_o;
  reg n9774_o;
  wire n9775_o;
  wire n9776_o;
  reg n9777_o;
  wire n9778_o;
  wire n9779_o;
  reg n9780_o;
  wire n9781_o;
  wire n9782_o;
  wire n9783_o;
  reg n9784_o;
  wire n9785_o;
  wire n9786_o;
  reg n9787_o;
  wire [31:0] n9810_o;
  wire [31:0] n9811_o;
  wire [20:0] n9812_o;
  wire [12:0] n9813_o;
  wire [31:0] n9814_o;
  assign ci_instr32_o = n9811_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:72:10  */
  assign imm20 = n9812_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:73:10  */
  assign imm12 = n9813_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:76:10  */
  assign illegal = n9747_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:77:10  */
  assign decoded = n9814_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:86:28  */
  assign n8990_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:87:28  */
  assign n8991_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:88:28  */
  assign n8992_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:89:28  */
  assign n8993_o = ci_instr16_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:90:28  */
  assign n8994_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:91:28  */
  assign n8995_o = ci_instr16_i[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:92:28  */
  assign n8996_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:93:28  */
  assign n8997_o = ci_instr16_i[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:94:28  */
  assign n8998_o = ci_instr16_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:95:28  */
  assign n8999_o = ci_instr16_i[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9000_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9001_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9002_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9003_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9004_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9005_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9006_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9007_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9008_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:96:49  */
  assign n9009_o = ci_instr16_i[12]; // extract
  assign n9010_o = {n9000_o, n9001_o, n9002_o, n9003_o};
  assign n9011_o = {n9004_o, n9005_o, n9006_o, n9007_o};
  assign n9012_o = {n9008_o, n9009_o};
  assign n9013_o = {n9010_o, n9011_o, n9012_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:100:28  */
  assign n9015_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:101:28  */
  assign n9016_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:102:28  */
  assign n9017_o = ci_instr16_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:103:28  */
  assign n9018_o = ci_instr16_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:104:28  */
  assign n9019_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:105:28  */
  assign n9020_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:106:28  */
  assign n9021_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:107:49  */
  assign n9022_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:107:49  */
  assign n9023_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:107:49  */
  assign n9024_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:107:49  */
  assign n9025_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:107:49  */
  assign n9026_o = ci_instr16_i[12]; // extract
  assign n9027_o = {n9022_o, n9023_o, n9024_o, n9025_o};
  assign n9028_o = {n9027_o, n9026_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:22  */
  assign n9030_o = ci_instr16_i[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:26  */
  assign n9031_o = ci_instr16_i[15:13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:128:89  */
  assign n9034_o = ci_instr16_i[4:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:128:75  */
  assign n9036_o = {2'b01, n9034_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:133:82  */
  assign n9043_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:134:82  */
  assign n9045_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:135:82  */
  assign n9047_o = ci_instr16_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:136:82  */
  assign n9049_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:137:82  */
  assign n9051_o = ci_instr16_i[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:138:82  */
  assign n9053_o = ci_instr16_i[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:139:82  */
  assign n9055_o = ci_instr16_i[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:140:82  */
  assign n9057_o = ci_instr16_i[10]; // extract
  assign n9058_o = n9038_o[11:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:141:29  */
  assign n9059_o = ci_instr16_i[12:5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:141:43  */
  assign n9061_o = n9059_o == 8'b00000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:141:13  */
  assign n9064_o = n9061_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:124:11  */
  assign n9066_o = n9031_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:149:82  */
  assign n9069_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:150:82  */
  assign n9070_o = ci_instr16_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:151:82  */
  assign n9071_o = ci_instr16_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:152:82  */
  assign n9072_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:153:82  */
  assign n9073_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:156:89  */
  assign n9076_o = ci_instr16_i[9:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:156:75  */
  assign n9078_o = {2'b01, n9076_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:157:89  */
  assign n9079_o = ci_instr16_i[4:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:157:75  */
  assign n9081_o = {2'b01, n9079_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:145:11  */
  assign n9083_o = n9031_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:163:82  */
  assign n9086_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:164:82  */
  assign n9087_o = ci_instr16_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:165:82  */
  assign n9088_o = ci_instr16_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:166:82  */
  assign n9089_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:167:82  */
  assign n9090_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:170:89  */
  assign n9093_o = ci_instr16_i[9:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:170:75  */
  assign n9095_o = {2'b01, n9093_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:171:89  */
  assign n9096_o = ci_instr16_i[4:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:171:75  */
  assign n9098_o = {2'b01, n9096_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:159:11  */
  assign n9100_o = n9031_o == 3'b110;
  assign n9101_o = {n9100_o, n9083_o, n9066_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9104_o = 1'b0;
      3'b010: n9104_o = 1'b0;
      3'b001: n9104_o = n9064_o;
      default: n9104_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9106_o = 7'b0100011;
      3'b010: n9106_o = 7'b0000011;
      3'b001: n9106_o = 7'b0010011;
      default: n9106_o = 7'b0000000;
    endcase
  assign n9107_o = n9036_o[1:0]; // extract
  assign n9108_o = n9081_o[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9110_o = 2'b00;
      3'b010: n9110_o = n9108_o;
      3'b001: n9110_o = n9107_o;
      default: n9110_o = 2'b00;
    endcase
  assign n9111_o = n9036_o[2]; // extract
  assign n9112_o = n9081_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9114_o = n9086_o;
      3'b010: n9114_o = n9112_o;
      3'b001: n9114_o = n9111_o;
      default: n9114_o = 1'b0;
    endcase
  assign n9115_o = n9036_o[3]; // extract
  assign n9116_o = n9081_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9118_o = n9087_o;
      3'b010: n9118_o = n9116_o;
      3'b001: n9118_o = n9115_o;
      default: n9118_o = 1'b0;
    endcase
  assign n9119_o = n9036_o[4]; // extract
  assign n9120_o = n9081_o[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9122_o = n9088_o;
      3'b010: n9122_o = n9120_o;
      3'b001: n9122_o = n9119_o;
      default: n9122_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9124_o = 3'b010;
      3'b010: n9124_o = 3'b010;
      3'b001: n9124_o = 3'b000;
      default: n9124_o = 3'b000;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9126_o = n9095_o;
      3'b010: n9126_o = n9078_o;
      3'b001: n9126_o = 5'b00010;
      default: n9126_o = 5'b00000;
    endcase
  assign n9127_o = n9068_o[0]; // extract
  assign n9128_o = n9098_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9130_o = n9128_o;
      3'b010: n9130_o = n9127_o;
      3'b001: n9130_o = 1'b0;
      default: n9130_o = 1'b0;
    endcase
  assign n9131_o = n9068_o[1]; // extract
  assign n9132_o = n9098_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9134_o = n9132_o;
      3'b010: n9134_o = n9131_o;
      3'b001: n9134_o = 1'b0;
      default: n9134_o = 1'b0;
    endcase
  assign n9135_o = n9098_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9137_o = n9135_o;
      3'b010: n9137_o = n9069_o;
      3'b001: n9137_o = n9043_o;
      default: n9137_o = 1'b0;
    endcase
  assign n9138_o = n9098_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9140_o = n9138_o;
      3'b010: n9140_o = n9070_o;
      3'b001: n9140_o = n9045_o;
      default: n9140_o = 1'b0;
    endcase
  assign n9141_o = n9098_o[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9143_o = n9141_o;
      3'b010: n9143_o = n9071_o;
      3'b001: n9143_o = n9047_o;
      default: n9143_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9145_o = n9089_o;
      3'b010: n9145_o = n9072_o;
      3'b001: n9145_o = n9049_o;
      default: n9145_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9147_o = n9090_o;
      3'b010: n9147_o = n9073_o;
      3'b001: n9147_o = n9051_o;
      default: n9147_o = 1'b0;
    endcase
  assign n9148_o = n9074_o[0]; // extract
  assign n9149_o = n9091_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9151_o = n9149_o;
      3'b010: n9151_o = n9148_o;
      3'b001: n9151_o = n9053_o;
      default: n9151_o = 1'b0;
    endcase
  assign n9152_o = n9074_o[1]; // extract
  assign n9153_o = n9091_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9155_o = n9153_o;
      3'b010: n9155_o = n9152_o;
      3'b001: n9155_o = n9055_o;
      default: n9155_o = 1'b0;
    endcase
  assign n9156_o = n9074_o[2]; // extract
  assign n9157_o = n9091_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9159_o = n9157_o;
      3'b010: n9159_o = n9156_o;
      3'b001: n9159_o = n9057_o;
      default: n9159_o = 1'b0;
    endcase
  assign n9160_o = n9074_o[4:3]; // extract
  assign n9161_o = n9091_o[4:3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:122:9  */
  always @*
    case (n9101_o)
      3'b100: n9163_o = n9161_o;
      3'b010: n9163_o = n9160_o;
      3'b001: n9163_o = n9058_o;
      default: n9163_o = 2'b00;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:121:7  */
  assign n9165_o = n9030_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:26  */
  assign n9166_o = ci_instr16_i[15:13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:184:29  */
  assign n9167_o = ci_instr16_i[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:184:13  */
  assign n9170_o = n9167_o ? 5'b00000 : 5'b00001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:190:75  */
  assign n9172_o = imm20[19:12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:191:75  */
  assign n9173_o = imm20[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:192:75  */
  assign n9174_o = imm20[10:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:193:75  */
  assign n9175_o = imm20[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:182:11  */
  assign n9177_o = n9166_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:182:22  */
  assign n9179_o = n9166_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:182:22  */
  assign n9180_o = n9177_o | n9179_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:197:29  */
  assign n9181_o = ci_instr16_i[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:197:47  */
  assign n9182_o = ~n9181_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:197:13  */
  assign n9185_o = n9182_o ? 3'b000 : 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:203:89  */
  assign n9187_o = ci_instr16_i[9:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:203:75  */
  assign n9189_o = {2'b01, n9187_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:205:75  */
  assign n9191_o = imm12[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:206:75  */
  assign n9192_o = imm12[4:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:207:75  */
  assign n9193_o = imm12[10:5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:208:75  */
  assign n9194_o = imm12[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:195:11  */
  assign n9196_o = n9166_o == 3'b110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:195:22  */
  assign n9198_o = n9166_o == 3'b111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:195:22  */
  assign n9199_o = n9196_o | n9198_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:215:82  */
  assign n9201_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9202_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9203_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9204_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9205_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9206_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9207_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9208_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9209_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9210_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9211_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9212_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:216:93  */
  assign n9213_o = ci_instr16_i[12]; // extract
  assign n9214_o = {n9202_o, n9203_o, n9204_o, n9205_o};
  assign n9215_o = {n9206_o, n9207_o, n9208_o, n9209_o};
  assign n9216_o = {n9210_o, n9211_o, n9212_o, n9213_o};
  assign n9217_o = {n9214_o, n9215_o, n9216_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:217:82  */
  assign n9218_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:218:82  */
  assign n9220_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:219:82  */
  assign n9222_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:220:82  */
  assign n9224_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:221:82  */
  assign n9226_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:222:82  */
  assign n9228_o = ci_instr16_i[12]; // extract
  assign n9229_o = n9217_o[11:6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:210:11  */
  assign n9231_o = n9166_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:226:29  */
  assign n9232_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:226:66  */
  assign n9234_o = n9232_o == 5'b00010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9238_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9239_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9240_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9241_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9242_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9243_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9244_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9245_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9246_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9247_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9248_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:232:95  */
  assign n9249_o = ci_instr16_i[12]; // extract
  assign n9250_o = {n9238_o, n9239_o, n9240_o, n9241_o};
  assign n9251_o = {n9242_o, n9243_o, n9244_o, n9245_o};
  assign n9252_o = {n9246_o, n9247_o, n9248_o, n9249_o};
  assign n9253_o = {n9250_o, n9251_o, n9252_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:237:84  */
  assign n9262_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:238:84  */
  assign n9264_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:239:84  */
  assign n9266_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:240:84  */
  assign n9268_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:241:84  */
  assign n9270_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:242:84  */
  assign n9272_o = ci_instr16_i[12]; // extract
  assign n9273_o = n9253_o[11:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:245:84  */
  assign n9275_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9276_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9277_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9278_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9279_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9280_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9281_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9282_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9283_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9284_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9285_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9286_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9287_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9288_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9289_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9290_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9291_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9292_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9293_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9294_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:246:95  */
  assign n9295_o = ci_instr16_i[12]; // extract
  assign n9296_o = {n9276_o, n9277_o, n9278_o, n9279_o};
  assign n9297_o = {n9280_o, n9281_o, n9282_o, n9283_o};
  assign n9298_o = {n9284_o, n9285_o, n9286_o, n9287_o};
  assign n9299_o = {n9288_o, n9289_o, n9290_o, n9291_o};
  assign n9300_o = {n9292_o, n9293_o, n9294_o, n9295_o};
  assign n9301_o = {n9296_o, n9297_o, n9298_o, n9299_o};
  assign n9302_o = {n9301_o, n9300_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:247:84  */
  assign n9303_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:248:84  */
  assign n9305_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:249:84  */
  assign n9307_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:250:84  */
  assign n9309_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:251:84  */
  assign n9311_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:252:84  */
  assign n9313_o = ci_instr16_i[12]; // extract
  assign n9314_o = n9302_o[19:6]; // extract
  assign n9315_o = {n9314_o, n9313_o, n9311_o, n9309_o, n9307_o, n9305_o, n9303_o, n9275_o, 7'b0110111};
  assign n9316_o = {n9273_o, n9272_o, n9270_o, n9268_o, n9266_o, n9264_o, n9262_o, 1'b0, 1'b0, 1'b0, 1'b0, 5'b00010, 3'b000, 5'b00010, 7'b0010011};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:226:13  */
  assign n9317_o = n9234_o ? n9316_o : n9315_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:254:29  */
  assign n9318_o = ci_instr16_i[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:254:42  */
  assign n9320_o = n9318_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:254:70  */
  assign n9321_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:254:75  */
  assign n9322_o = ~n9321_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:254:53  */
  assign n9323_o = n9322_o & n9320_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:254:13  */
  assign n9326_o = n9323_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:224:11  */
  assign n9328_o = n9166_o == 3'b011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:262:82  */
  assign n9329_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:263:82  */
  assign n9330_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9331_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9332_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9333_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9334_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9335_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9336_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9337_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9338_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9339_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9340_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9341_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:264:93  */
  assign n9342_o = ci_instr16_i[12]; // extract
  assign n9343_o = {n9331_o, n9332_o, n9333_o, n9334_o};
  assign n9344_o = {n9335_o, n9336_o, n9337_o, n9338_o};
  assign n9345_o = {n9339_o, n9340_o, n9341_o, n9342_o};
  assign n9346_o = {n9343_o, n9344_o, n9345_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:265:82  */
  assign n9347_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:266:82  */
  assign n9349_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:267:82  */
  assign n9351_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:268:82  */
  assign n9353_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:269:82  */
  assign n9355_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:270:82  */
  assign n9357_o = ci_instr16_i[12]; // extract
  assign n9358_o = n9346_o[11:6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:258:11  */
  assign n9360_o = n9166_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:274:83  */
  assign n9361_o = ci_instr16_i[9:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:274:69  */
  assign n9363_o = {2'b01, n9361_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:275:83  */
  assign n9364_o = ci_instr16_i[9:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:275:69  */
  assign n9366_o = {2'b01, n9364_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:276:83  */
  assign n9367_o = ci_instr16_i[4:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:276:69  */
  assign n9369_o = {2'b01, n9367_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:30  */
  assign n9370_o = ci_instr16_i[11:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:279:33  */
  assign n9371_o = ci_instr16_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:279:38  */
  assign n9372_o = ~n9371_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:279:17  */
  assign n9375_o = n9372_o ? 7'b0000000 : 7'b0100000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:286:86  */
  assign n9377_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:287:86  */
  assign n9378_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:288:86  */
  assign n9379_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:289:86  */
  assign n9380_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:290:86  */
  assign n9381_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:291:33  */
  assign n9382_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:291:17  */
  assign n9385_o = n9382_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:278:15  */
  assign n9387_o = n9370_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:278:25  */
  assign n9389_o = n9370_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:278:25  */
  assign n9390_o = n9387_o | n9389_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9392_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9393_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9394_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9395_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9396_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9397_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9398_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9399_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9400_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9401_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9402_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:297:97  */
  assign n9403_o = ci_instr16_i[12]; // extract
  assign n9404_o = {n9392_o, n9393_o, n9394_o, n9395_o};
  assign n9405_o = {n9396_o, n9397_o, n9398_o, n9399_o};
  assign n9406_o = {n9400_o, n9401_o, n9402_o, n9403_o};
  assign n9407_o = {n9404_o, n9405_o, n9406_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:298:86  */
  assign n9408_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:299:86  */
  assign n9410_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:300:86  */
  assign n9412_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:301:86  */
  assign n9414_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:302:86  */
  assign n9416_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:303:86  */
  assign n9418_o = ci_instr16_i[12]; // extract
  assign n9419_o = n9407_o[11:6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:294:15  */
  assign n9421_o = n9370_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:306:34  */
  assign n9423_o = ci_instr16_i[6:5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:307:19  */
  assign n9426_o = n9423_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:310:19  */
  assign n9430_o = n9423_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:313:19  */
  assign n9434_o = n9423_o == 2'b10;
  assign n9436_o = {n9434_o, n9430_o, n9426_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:306:17  */
  always @*
    case (n9436_o)
      3'b100: n9437_o = 3'b110;
      3'b010: n9437_o = 3'b100;
      3'b001: n9437_o = 3'b000;
      default: n9437_o = 3'b111;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:306:17  */
  always @*
    case (n9436_o)
      3'b100: n9438_o = 7'b0000000;
      3'b010: n9438_o = 7'b0000000;
      3'b001: n9438_o = 7'b0100000;
      default: n9438_o = 7'b0000000;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:320:33  */
  assign n9439_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:320:17  */
  assign n9442_o = n9439_o ? 1'b1 : 1'b0;
  assign n9443_o = {n9421_o, n9390_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9445_o = 1'b0;
      2'b01: n9445_o = n9385_o;
      default: n9445_o = n9442_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9446_o = 7'b0010011;
      2'b01: n9446_o = 7'b0010011;
      default: n9446_o = 7'b0110011;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9447_o = 3'b111;
      2'b01: n9447_o = 3'b101;
      default: n9447_o = n9437_o;
    endcase
  assign n9448_o = n9369_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9449_o = n9408_o;
      2'b01: n9449_o = n9377_o;
      default: n9449_o = n9448_o;
    endcase
  assign n9450_o = n9369_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9451_o = n9410_o;
      2'b01: n9451_o = n9378_o;
      default: n9451_o = n9450_o;
    endcase
  assign n9452_o = n9369_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9453_o = n9412_o;
      2'b01: n9453_o = n9379_o;
      default: n9453_o = n9452_o;
    endcase
  assign n9454_o = n9369_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9455_o = n9414_o;
      2'b01: n9455_o = n9380_o;
      default: n9455_o = n9454_o;
    endcase
  assign n9456_o = n9369_o[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9457_o = n9416_o;
      2'b01: n9457_o = n9381_o;
      default: n9457_o = n9456_o;
    endcase
  assign n9458_o = n9375_o[0]; // extract
  assign n9459_o = n9438_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9460_o = n9418_o;
      2'b01: n9460_o = n9458_o;
      default: n9460_o = n9459_o;
    endcase
  assign n9461_o = n9375_o[6:1]; // extract
  assign n9462_o = n9438_o[6:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:277:13  */
  always @*
    case (n9443_o)
      2'b10: n9463_o = n9419_o;
      2'b01: n9463_o = n9461_o;
      default: n9463_o = n9462_o;
    endcase
  assign n9468_o = {n9360_o, n9328_o, n9231_o, n9199_o, n9180_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9470_o = 1'b0;
      5'b01000: n9470_o = n9326_o;
      5'b00100: n9470_o = 1'b0;
      5'b00010: n9470_o = 1'b0;
      5'b00001: n9470_o = 1'b0;
      default: n9470_o = n9445_o;
    endcase
  assign n9471_o = n9317_o[6:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9472_o = 7'b0010011;
      5'b01000: n9472_o = n9471_o;
      5'b00100: n9472_o = 7'b0010011;
      5'b00010: n9472_o = 7'b1100011;
      5'b00001: n9472_o = 7'b1101111;
      default: n9472_o = n9446_o;
    endcase
  assign n9473_o = n9170_o[0]; // extract
  assign n9474_o = n9201_o[0]; // extract
  assign n9475_o = n9317_o[7]; // extract
  assign n9476_o = n9330_o[0]; // extract
  assign n9477_o = n9363_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9478_o = n9476_o;
      5'b01000: n9478_o = n9475_o;
      5'b00100: n9478_o = n9474_o;
      5'b00010: n9478_o = n9191_o;
      5'b00001: n9478_o = n9473_o;
      default: n9478_o = n9477_o;
    endcase
  assign n9479_o = n9170_o[4:1]; // extract
  assign n9480_o = n9201_o[4:1]; // extract
  assign n9481_o = n9317_o[11:8]; // extract
  assign n9482_o = n9330_o[4:1]; // extract
  assign n9483_o = n9363_o[4:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9484_o = n9482_o;
      5'b01000: n9484_o = n9481_o;
      5'b00100: n9484_o = n9480_o;
      5'b00010: n9484_o = n9192_o;
      5'b00001: n9484_o = n9479_o;
      default: n9484_o = n9483_o;
    endcase
  assign n9485_o = n9172_o[2:0]; // extract
  assign n9486_o = n9317_o[14:12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9487_o = 3'b000;
      5'b01000: n9487_o = n9486_o;
      5'b00100: n9487_o = 3'b000;
      5'b00010: n9487_o = n9185_o;
      5'b00001: n9487_o = n9485_o;
      default: n9487_o = n9447_o;
    endcase
  assign n9488_o = n9172_o[7:3]; // extract
  assign n9489_o = n9317_o[19:15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9490_o = n9329_o;
      5'b01000: n9490_o = n9489_o;
      5'b00100: n9490_o = 5'b00000;
      5'b00010: n9490_o = n9189_o;
      5'b00001: n9490_o = n9488_o;
      default: n9490_o = n9366_o;
    endcase
  assign n9491_o = n9190_o[0]; // extract
  assign n9492_o = n9317_o[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9493_o = n9347_o;
      5'b01000: n9493_o = n9492_o;
      5'b00100: n9493_o = n9218_o;
      5'b00010: n9493_o = n9491_o;
      5'b00001: n9493_o = n9173_o;
      default: n9493_o = n9449_o;
    endcase
  assign n9494_o = n9174_o[0]; // extract
  assign n9495_o = n9190_o[1]; // extract
  assign n9496_o = n9317_o[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9497_o = n9349_o;
      5'b01000: n9497_o = n9496_o;
      5'b00100: n9497_o = n9220_o;
      5'b00010: n9497_o = n9495_o;
      5'b00001: n9497_o = n9494_o;
      default: n9497_o = n9451_o;
    endcase
  assign n9498_o = n9174_o[1]; // extract
  assign n9499_o = n9190_o[2]; // extract
  assign n9500_o = n9317_o[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9501_o = n9351_o;
      5'b01000: n9501_o = n9500_o;
      5'b00100: n9501_o = n9222_o;
      5'b00010: n9501_o = n9499_o;
      5'b00001: n9501_o = n9498_o;
      default: n9501_o = n9453_o;
    endcase
  assign n9502_o = n9174_o[2]; // extract
  assign n9503_o = n9190_o[3]; // extract
  assign n9504_o = n9317_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9505_o = n9353_o;
      5'b01000: n9505_o = n9504_o;
      5'b00100: n9505_o = n9224_o;
      5'b00010: n9505_o = n9503_o;
      5'b00001: n9505_o = n9502_o;
      default: n9505_o = n9455_o;
    endcase
  assign n9506_o = n9174_o[3]; // extract
  assign n9507_o = n9190_o[4]; // extract
  assign n9508_o = n9317_o[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9509_o = n9355_o;
      5'b01000: n9509_o = n9508_o;
      5'b00100: n9509_o = n9226_o;
      5'b00010: n9509_o = n9507_o;
      5'b00001: n9509_o = n9506_o;
      default: n9509_o = n9457_o;
    endcase
  assign n9510_o = n9174_o[4]; // extract
  assign n9511_o = n9193_o[0]; // extract
  assign n9512_o = n9317_o[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9513_o = n9357_o;
      5'b01000: n9513_o = n9512_o;
      5'b00100: n9513_o = n9228_o;
      5'b00010: n9513_o = n9511_o;
      5'b00001: n9513_o = n9510_o;
      default: n9513_o = n9460_o;
    endcase
  assign n9514_o = n9174_o[9:5]; // extract
  assign n9515_o = n9193_o[5:1]; // extract
  assign n9516_o = n9229_o[4:0]; // extract
  assign n9517_o = n9317_o[30:26]; // extract
  assign n9518_o = n9358_o[4:0]; // extract
  assign n9519_o = n9463_o[4:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9520_o = n9518_o;
      5'b01000: n9520_o = n9517_o;
      5'b00100: n9520_o = n9516_o;
      5'b00010: n9520_o = n9515_o;
      5'b00001: n9520_o = n9514_o;
      default: n9520_o = n9519_o;
    endcase
  assign n9521_o = n9229_o[5]; // extract
  assign n9522_o = n9317_o[31]; // extract
  assign n9523_o = n9358_o[5]; // extract
  assign n9524_o = n9463_o[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:181:9  */
  always @*
    case (n9468_o)
      5'b10000: n9525_o = n9523_o;
      5'b01000: n9525_o = n9522_o;
      5'b00100: n9525_o = n9521_o;
      5'b00010: n9525_o = n9194_o;
      5'b00001: n9525_o = n9175_o;
      default: n9525_o = n9524_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:179:7  */
  assign n9527_o = n9030_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:26  */
  assign n9528_o = ci_instr16_i[15:13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:333:82  */
  assign n9529_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:334:82  */
  assign n9530_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:337:82  */
  assign n9533_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:338:82  */
  assign n9534_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:339:82  */
  assign n9535_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:340:82  */
  assign n9536_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:341:82  */
  assign n9537_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:342:29  */
  assign n9538_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:342:13  */
  assign n9541_o = n9538_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:330:11  */
  assign n9543_o = n9528_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:350:82  */
  assign n9545_o = ci_instr16_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:351:82  */
  assign n9546_o = ci_instr16_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:352:82  */
  assign n9547_o = ci_instr16_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:353:82  */
  assign n9548_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:354:82  */
  assign n9549_o = ci_instr16_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:355:82  */
  assign n9550_o = ci_instr16_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:359:82  */
  assign n9553_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:360:29  */
  assign n9554_o = ci_instr16_i[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:361:29  */
  assign n9555_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:361:66  */
  assign n9557_o = n9555_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:360:54  */
  assign n9558_o = n9554_o | n9557_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:360:13  */
  assign n9561_o = n9558_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:346:11  */
  assign n9563_o = n9528_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:346:22  */
  assign n9565_o = n9528_o == 3'b011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:346:22  */
  assign n9566_o = n9563_o | n9565_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:369:82  */
  assign n9568_o = ci_instr16_i[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:370:82  */
  assign n9569_o = ci_instr16_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:371:82  */
  assign n9570_o = ci_instr16_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:372:82  */
  assign n9571_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:373:82  */
  assign n9572_o = ci_instr16_i[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:374:82  */
  assign n9573_o = ci_instr16_i[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:378:82  */
  assign n9576_o = ci_instr16_i[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:379:29  */
  assign n9577_o = ci_instr16_i[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:379:13  */
  assign n9580_o = n9577_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:365:11  */
  assign n9582_o = n9528_o == 3'b110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:365:22  */
  assign n9584_o = n9528_o == 3'b111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:365:22  */
  assign n9585_o = n9582_o | n9584_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:385:29  */
  assign n9586_o = ci_instr16_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:385:34  */
  assign n9587_o = ~n9586_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:386:31  */
  assign n9588_o = ci_instr16_i[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:386:44  */
  assign n9590_o = n9588_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:388:86  */
  assign n9592_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:390:33  */
  assign n9594_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:390:72  */
  assign n9596_o = n9594_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:391:33  */
  assign n9597_o = ci_instr16_i[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:391:72  */
  assign n9599_o = n9597_o != 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:390:83  */
  assign n9600_o = n9596_o | n9599_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:390:17  */
  assign n9603_o = n9600_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:397:86  */
  assign n9605_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:399:86  */
  assign n9607_o = ci_instr16_i[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:400:33  */
  assign n9608_o = ci_instr16_i[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:400:72  */
  assign n9610_o = n9608_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:400:17  */
  assign n9613_o = n9610_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:386:15  */
  assign n9614_o = n9590_o ? n9603_o : n9613_o;
  assign n9615_o = {n9607_o, 5'b00000, 3'b000, n9605_o, 7'b0110011};
  assign n9616_o = {5'b00000, 7'b1100111};
  assign n9617_o = n9615_o[11:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:386:15  */
  assign n9618_o = n9590_o ? n9616_o : n9617_o;
  assign n9619_o = n9615_o[14:12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:386:15  */
  assign n9621_o = n9590_o ? 3'b000 : n9619_o;
  assign n9622_o = n9615_o[19:15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:386:15  */
  assign n9623_o = n9590_o ? n9592_o : n9622_o;
  assign n9624_o = n9615_o[24:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:386:15  */
  assign n9626_o = n9590_o ? 5'b00000 : n9624_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:405:31  */
  assign n9627_o = ci_instr16_i[6:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:405:44  */
  assign n9629_o = n9627_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:406:33  */
  assign n9630_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:406:47  */
  assign n9632_o = n9630_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:411:88  */
  assign n9635_o = ci_instr16_i[11:7]; // extract
  assign n9637_o = {5'b00001, 7'b1100111};
  assign n9638_o = n9637_o[6:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:406:17  */
  assign n9639_o = n9632_o ? 7'b1110011 : n9638_o;
  assign n9640_o = n9637_o[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:406:17  */
  assign n9642_o = n9632_o ? 5'b00000 : n9640_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:406:17  */
  assign n9644_o = n9632_o ? 5'b00000 : n9635_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:406:17  */
  assign n9646_o = n9632_o ? 12'b000000000001 : 12'b000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:417:86  */
  assign n9648_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:418:86  */
  assign n9649_o = ci_instr16_i[11:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:419:86  */
  assign n9650_o = ci_instr16_i[6:2]; // extract
  assign n9651_o = {n9650_o, n9649_o, 3'b000, n9648_o, 7'b0110011};
  assign n9652_o = {n9642_o, n9639_o};
  assign n9653_o = {n9646_o, n9644_o};
  assign n9654_o = n9651_o[11:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:405:15  */
  assign n9655_o = n9629_o ? n9652_o : n9654_o;
  assign n9656_o = n9651_o[14:12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:405:15  */
  assign n9658_o = n9629_o ? 3'b000 : n9656_o;
  assign n9659_o = n9651_o[24:15]; // extract
  assign n9660_o = n9653_o[9:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:405:15  */
  assign n9661_o = n9629_o ? n9660_o : n9659_o;
  assign n9662_o = n9653_o[16:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:405:15  */
  assign n9664_o = n9629_o ? n9662_o : 7'b0000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:385:13  */
  assign n9666_o = n9587_o ? n9614_o : 1'b0;
  assign n9667_o = {n9664_o, n9661_o, n9658_o, n9655_o};
  assign n9668_o = {n9626_o, n9623_o, n9621_o, n9618_o};
  assign n9669_o = n9667_o[24:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:385:13  */
  assign n9670_o = n9587_o ? n9668_o : n9669_o;
  assign n9671_o = n9667_o[31:25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:385:13  */
  assign n9673_o = n9587_o ? 7'b0000000 : n9671_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:383:11  */
  assign n9675_o = n9528_o == 3'b100;
  assign n9676_o = {n9675_o, n9585_o, n9566_o, n9543_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9678_o = n9666_o;
      4'b0100: n9678_o = n9580_o;
      4'b0010: n9678_o = n9561_o;
      4'b0001: n9678_o = n9541_o;
      default: n9678_o = 1'b1;
    endcase
  assign n9679_o = n9670_o[6:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9681_o = n9679_o;
      4'b0100: n9681_o = 7'b0100011;
      4'b0010: n9681_o = 7'b0000011;
      4'b0001: n9681_o = 7'b0010011;
      default: n9681_o = 7'b0000000;
    endcase
  assign n9682_o = n9530_o[1:0]; // extract
  assign n9683_o = n9553_o[1:0]; // extract
  assign n9684_o = n9670_o[8:7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9686_o = n9684_o;
      4'b0100: n9686_o = 2'b00;
      4'b0010: n9686_o = n9683_o;
      4'b0001: n9686_o = n9682_o;
      default: n9686_o = 2'b00;
    endcase
  assign n9687_o = n9530_o[2]; // extract
  assign n9688_o = n9553_o[2]; // extract
  assign n9689_o = n9670_o[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9691_o = n9689_o;
      4'b0100: n9691_o = n9568_o;
      4'b0010: n9691_o = n9688_o;
      4'b0001: n9691_o = n9687_o;
      default: n9691_o = 1'b0;
    endcase
  assign n9692_o = n9530_o[3]; // extract
  assign n9693_o = n9553_o[3]; // extract
  assign n9694_o = n9670_o[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9696_o = n9694_o;
      4'b0100: n9696_o = n9569_o;
      4'b0010: n9696_o = n9693_o;
      4'b0001: n9696_o = n9692_o;
      default: n9696_o = 1'b0;
    endcase
  assign n9697_o = n9530_o[4]; // extract
  assign n9698_o = n9553_o[4]; // extract
  assign n9699_o = n9670_o[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9701_o = n9699_o;
      4'b0100: n9701_o = n9570_o;
      4'b0010: n9701_o = n9698_o;
      4'b0001: n9701_o = n9697_o;
      default: n9701_o = 1'b0;
    endcase
  assign n9702_o = n9670_o[14:12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9704_o = n9702_o;
      4'b0100: n9704_o = 3'b010;
      4'b0010: n9704_o = 3'b010;
      4'b0001: n9704_o = 3'b001;
      default: n9704_o = 3'b000;
    endcase
  assign n9705_o = n9670_o[19:15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9707_o = n9705_o;
      4'b0100: n9707_o = 5'b00010;
      4'b0010: n9707_o = 5'b00010;
      4'b0001: n9707_o = n9529_o;
      default: n9707_o = 5'b00000;
    endcase
  assign n9708_o = n9544_o[0]; // extract
  assign n9709_o = n9576_o[0]; // extract
  assign n9710_o = n9670_o[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9712_o = n9710_o;
      4'b0100: n9712_o = n9709_o;
      4'b0010: n9712_o = n9708_o;
      4'b0001: n9712_o = n9533_o;
      default: n9712_o = 1'b0;
    endcase
  assign n9713_o = n9544_o[1]; // extract
  assign n9714_o = n9576_o[1]; // extract
  assign n9715_o = n9670_o[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9717_o = n9715_o;
      4'b0100: n9717_o = n9714_o;
      4'b0010: n9717_o = n9713_o;
      4'b0001: n9717_o = n9534_o;
      default: n9717_o = 1'b0;
    endcase
  assign n9718_o = n9576_o[2]; // extract
  assign n9719_o = n9670_o[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9721_o = n9719_o;
      4'b0100: n9721_o = n9718_o;
      4'b0010: n9721_o = n9545_o;
      4'b0001: n9721_o = n9535_o;
      default: n9721_o = 1'b0;
    endcase
  assign n9722_o = n9576_o[3]; // extract
  assign n9723_o = n9670_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9725_o = n9723_o;
      4'b0100: n9725_o = n9722_o;
      4'b0010: n9725_o = n9546_o;
      4'b0001: n9725_o = n9536_o;
      default: n9725_o = 1'b0;
    endcase
  assign n9726_o = n9576_o[4]; // extract
  assign n9727_o = n9670_o[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9729_o = n9727_o;
      4'b0100: n9729_o = n9726_o;
      4'b0010: n9729_o = n9547_o;
      4'b0001: n9729_o = n9537_o;
      default: n9729_o = 1'b0;
    endcase
  assign n9730_o = n9532_o[0]; // extract
  assign n9731_o = n9673_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9733_o = n9731_o;
      4'b0100: n9733_o = n9571_o;
      4'b0010: n9733_o = n9548_o;
      4'b0001: n9733_o = n9730_o;
      default: n9733_o = 1'b0;
    endcase
  assign n9734_o = n9532_o[1]; // extract
  assign n9735_o = n9673_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9737_o = n9735_o;
      4'b0100: n9737_o = n9572_o;
      4'b0010: n9737_o = n9549_o;
      4'b0001: n9737_o = n9734_o;
      default: n9737_o = 1'b0;
    endcase
  assign n9738_o = n9532_o[2]; // extract
  assign n9739_o = n9673_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9741_o = n9739_o;
      4'b0100: n9741_o = n9573_o;
      4'b0010: n9741_o = n9550_o;
      4'b0001: n9741_o = n9738_o;
      default: n9741_o = 1'b0;
    endcase
  assign n9742_o = n9532_o[6:3]; // extract
  assign n9743_o = n9673_o[6:3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:328:9  */
  always @*
    case (n9676_o)
      4'b1000: n9745_o = n9743_o;
      4'b0100: n9745_o = 4'b0000;
      4'b0010: n9745_o = 4'b0000;
      4'b0001: n9745_o = n9742_o;
      default: n9745_o = 4'b0000;
    endcase
  assign n9746_o = {n9527_o, n9165_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9747_o = n9470_o;
      2'b01: n9747_o = n9104_o;
      default: n9747_o = n9678_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9749_o = n9472_o;
      2'b01: n9749_o = n9106_o;
      default: n9749_o = n9681_o;
    endcase
  assign n9750_o = n9110_o[0]; // extract
  assign n9751_o = n9686_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9752_o = n9478_o;
      2'b01: n9752_o = n9750_o;
      default: n9752_o = n9751_o;
    endcase
  assign n9753_o = n9110_o[1]; // extract
  assign n9754_o = n9484_o[0]; // extract
  assign n9755_o = n9686_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9756_o = n9754_o;
      2'b01: n9756_o = n9753_o;
      default: n9756_o = n9755_o;
    endcase
  assign n9757_o = n9484_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9758_o = n9757_o;
      2'b01: n9758_o = n9114_o;
      default: n9758_o = n9691_o;
    endcase
  assign n9759_o = n9484_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9760_o = n9759_o;
      2'b01: n9760_o = n9118_o;
      default: n9760_o = n9696_o;
    endcase
  assign n9761_o = n9484_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9762_o = n9761_o;
      2'b01: n9762_o = n9122_o;
      default: n9762_o = n9701_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9763_o = n9487_o;
      2'b01: n9763_o = n9124_o;
      default: n9763_o = n9704_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9764_o = n9490_o;
      2'b01: n9764_o = n9126_o;
      default: n9764_o = n9707_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9765_o = n9493_o;
      2'b01: n9765_o = n9130_o;
      default: n9765_o = n9712_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9766_o = n9497_o;
      2'b01: n9766_o = n9134_o;
      default: n9766_o = n9717_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9767_o = n9501_o;
      2'b01: n9767_o = n9137_o;
      default: n9767_o = n9721_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9768_o = n9505_o;
      2'b01: n9768_o = n9140_o;
      default: n9768_o = n9725_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9769_o = n9509_o;
      2'b01: n9769_o = n9143_o;
      default: n9769_o = n9729_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9770_o = n9513_o;
      2'b01: n9770_o = n9145_o;
      default: n9770_o = n9733_o;
    endcase
  assign n9771_o = n9520_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9772_o = n9771_o;
      2'b01: n9772_o = n9147_o;
      default: n9772_o = n9737_o;
    endcase
  assign n9773_o = n9520_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9774_o = n9773_o;
      2'b01: n9774_o = n9151_o;
      default: n9774_o = n9741_o;
    endcase
  assign n9775_o = n9520_o[2]; // extract
  assign n9776_o = n9745_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9777_o = n9775_o;
      2'b01: n9777_o = n9155_o;
      default: n9777_o = n9776_o;
    endcase
  assign n9778_o = n9520_o[3]; // extract
  assign n9779_o = n9745_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9780_o = n9778_o;
      2'b01: n9780_o = n9159_o;
      default: n9780_o = n9779_o;
    endcase
  assign n9781_o = n9163_o[0]; // extract
  assign n9782_o = n9520_o[4]; // extract
  assign n9783_o = n9745_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9784_o = n9782_o;
      2'b01: n9784_o = n9781_o;
      default: n9784_o = n9783_o;
    endcase
  assign n9785_o = n9163_o[1]; // extract
  assign n9786_o = n9745_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:119:5  */
  always @*
    case (n9746_o)
      2'b10: n9787_o = n9525_o;
      2'b01: n9787_o = n9785_o;
      default: n9787_o = n9786_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:433:28  */
  assign n9810_o = {16'b0000000000000000, ci_instr16_i};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_decompressor.vhd:433:44  */
  assign n9811_o = illegal ? n9810_o : decoded;
  assign n9812_o = {n9013_o, n8999_o, n8998_o, n8997_o, n8996_o, n8995_o, n8994_o, n8993_o, n8992_o, n8991_o, n8990_o, 1'b0};
  assign n9813_o = {n9028_o, n9021_o, n9020_o, n9019_o, n9018_o, n9017_o, n9016_o, n9015_o, 1'b0};
  assign n9814_o = {n9787_o, n9784_o, n9780_o, n9777_o, n9774_o, n9772_o, n9770_o, n9769_o, n9768_o, n9767_o, n9766_o, n9765_o, n9764_o, n9763_o, n9762_o, n9760_o, n9758_o, n9756_o, n9752_o, n9749_o};
endmodule

module neorv32_fifo_2_17_29e2dcfbb16f63bb0254df7585a15bb6fb5e927d
  (input  clk_i,
   input  rstn_i,
   input  clear_i,
   input  [16:0] wdata_i,
   input  we_i,
   input  re_i,
   output half_o,
   output free_o,
   output [16:0] rdata_o,
   output avail_o);
  wire we;
  wire re;
  wire [1:0] w_pnt;
  wire [1:0] r_pnt;
  wire [1:0] w_nxt;
  wire [1:0] r_nxt;
  wire [1:0] r_pnt_ff;
  wire match;
  wire empty;
  wire full;
  wire half;
  wire free;
  wire avail;
  wire [1:0] diff;
  wire n8909_o;
  wire n8910_o;
  wire n8912_o;
  wire n8913_o;
  wire n8915_o;
  wire [1:0] n8925_o;
  wire [1:0] n8927_o;
  wire [1:0] n8928_o;
  wire [1:0] n8930_o;
  wire [1:0] n8932_o;
  wire [1:0] n8933_o;
  wire n8935_o;
  wire n8936_o;
  wire n8937_o;
  wire n8938_o;
  wire n8941_o;
  wire n8942_o;
  wire n8943_o;
  wire n8944_o;
  wire n8945_o;
  wire n8948_o;
  wire n8949_o;
  wire n8950_o;
  wire n8951_o;
  wire n8952_o;
  wire [1:0] n8954_o;
  wire n8955_o;
  wire n8956_o;
  wire n8957_o;
  wire n8958_o;
  wire n8961_o;
  wire n8974_o;
  reg [1:0] n8983_q;
  reg [1:0] n8984_q;
  reg [1:0] n8985_q;
  wire [16:0] n8986_data; // mem_rd
  assign half_o = half; //(module output)
  assign free_o = free; //(module output)
  assign rdata_o = n8986_data; //(module output)
  assign avail_o = avail; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:77:10  */
  assign we = n8912_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:77:17  */
  assign re = n8909_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:78:10  */
  assign w_pnt = n8983_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:78:17  */
  assign r_pnt = n8984_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:79:10  */
  assign w_nxt = n8925_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:79:17  */
  assign r_nxt = n8930_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:82:10  */
  assign r_pnt_ff = n8985_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:85:10  */
  assign match = n8938_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:85:17  */
  assign empty = n8952_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:85:24  */
  assign full = n8945_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:85:30  */
  assign half = n8956_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:85:36  */
  assign free = n8957_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:85:42  */
  assign avail = n8958_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:88:10  */
  assign diff = n8954_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:94:14  */
  assign n8909_o = 1'b1 ? re_i : n8910_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:94:50  */
  assign n8910_o = re_i & avail;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:95:14  */
  assign n8912_o = 1'b1 ? we_i : n8913_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:95:50  */
  assign n8913_o = we_i & free;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:102:16  */
  assign n8915_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:112:28  */
  assign n8925_o = clear_i ? 2'b00 : n8928_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:112:88  */
  assign n8927_o = w_pnt + 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:112:49  */
  assign n8928_o = we ? n8927_o : w_pnt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:113:28  */
  assign n8930_o = clear_i ? 2'b00 : n8933_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:113:88  */
  assign n8932_o = r_pnt + 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:113:49  */
  assign n8933_o = re ? n8932_o : r_pnt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:122:29  */
  assign n8935_o = r_pnt[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:122:60  */
  assign n8936_o = w_pnt[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:122:53  */
  assign n8937_o = n8935_o == n8936_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:122:18  */
  assign n8938_o = n8937_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:123:29  */
  assign n8941_o = r_pnt[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:123:50  */
  assign n8942_o = w_pnt[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:123:42  */
  assign n8943_o = n8941_o != n8942_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:123:64  */
  assign n8944_o = match & n8943_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:123:18  */
  assign n8945_o = n8944_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:124:29  */
  assign n8948_o = r_pnt[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:124:50  */
  assign n8949_o = w_pnt[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:124:43  */
  assign n8950_o = n8948_o == n8949_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:124:64  */
  assign n8951_o = match & n8950_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:124:18  */
  assign n8952_o = n8951_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:125:48  */
  assign n8954_o = w_pnt - r_pnt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:126:18  */
  assign n8955_o = diff[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:126:32  */
  assign n8956_o = n8955_o | full;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:138:12  */
  assign n8957_o = ~full;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:139:12  */
  assign n8958_o = ~empty;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:205:47  */
  assign n8961_o = w_pnt[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:234:55  */
  assign n8974_o = r_pnt_ff[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:105:5  */
  always @(posedge clk_i or posedge n8915_o)
    if (n8915_o)
      n8983_q <= 2'b00;
    else
      n8983_q <= w_nxt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:105:5  */
  always @(posedge clk_i or posedge n8915_o)
    if (n8915_o)
      n8984_q <= 2'b00;
    else
      n8984_q <= r_nxt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:230:9  */
  always @(posedge clk_i)
    n8985_q <= r_nxt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:234:27  */
  reg [16:0] fifo_mem[1:0] ; // memory
  assign n8986_data = fifo_mem[n8974_o];
  always @(posedge clk_i)
    if (we)
      fifo_mem[n8961_o] <= wdata_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:234:27  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_fifo.vhd:205:22  */
endmodule

module neorv32_bus_switch_1489f923c4dca729178b3e3233458550d8dddf29
  (input  clk_i,
   input  rstn_i,
   input  [31:0] a_req_i_addr,
   input  [31:0] a_req_i_data,
   input  [3:0] a_req_i_ben,
   input  a_req_i_stb,
   input  a_req_i_rw,
   input  a_req_i_src,
   input  a_req_i_priv,
   input  a_req_i_rvso,
   input  a_req_i_fence,
   input  [31:0] b_req_i_addr,
   input  [31:0] b_req_i_data,
   input  [3:0] b_req_i_ben,
   input  b_req_i_stb,
   input  b_req_i_rw,
   input  b_req_i_src,
   input  b_req_i_priv,
   input  b_req_i_rvso,
   input  b_req_i_fence,
   input  [31:0] x_rsp_i_data,
   input  x_rsp_i_ack,
   input  x_rsp_i_err,
   output [31:0] a_rsp_o_data,
   output a_rsp_o_ack,
   output a_rsp_o_err,
   output [31:0] b_rsp_o_data,
   output b_rsp_o_ack,
   output b_rsp_o_err,
   output [31:0] x_req_o_addr,
   output [31:0] x_req_o_data,
   output [3:0] x_req_o_ben,
   output x_req_o_stb,
   output x_req_o_rw,
   output x_req_o_src,
   output x_req_o_priv,
   output x_req_o_rvso,
   output x_req_o_fence);
  wire [73:0] n8733_o;
  wire [31:0] n8735_o;
  wire n8736_o;
  wire n8737_o;
  wire [73:0] n8738_o;
  wire [31:0] n8740_o;
  wire n8741_o;
  wire n8742_o;
  wire [31:0] n8744_o;
  wire [31:0] n8745_o;
  wire [3:0] n8746_o;
  wire n8747_o;
  wire n8748_o;
  wire n8749_o;
  wire n8750_o;
  wire n8751_o;
  wire n8752_o;
  wire [33:0] n8753_o;
  wire [7:0] arbiter;
  wire n8755_o;
  wire [1:0] n8760_o;
  wire n8761_o;
  wire n8762_o;
  wire n8763_o;
  wire n8764_o;
  wire n8765_o;
  wire n8766_o;
  wire n8767_o;
  wire n8768_o;
  wire n8769_o;
  wire n8770_o;
  wire n8771_o;
  wire n8772_o;
  wire [1:0] n8773_o;
  wire [1:0] n8778_o;
  wire [1:0] n8783_o;
  wire [1:0] n8786_o;
  wire n8788_o;
  wire n8789_o;
  wire n8790_o;
  wire [1:0] n8791_o;
  wire n8793_o;
  wire n8795_o;
  wire n8796_o;
  wire n8797_o;
  wire [1:0] n8798_o;
  wire n8800_o;
  wire n8801_o;
  wire n8802_o;
  wire n8803_o;
  wire n8807_o;
  wire n8808_o;
  wire n8809_o;
  wire [1:0] n8813_o;
  wire [1:0] n8814_o;
  wire [1:0] n8815_o;
  wire [1:0] n8816_o;
  wire [1:0] n8817_o;
  wire [1:0] n8818_o;
  wire [1:0] n8819_o;
  wire [1:0] n8820_o;
  reg [1:0] n8821_o;
  wire n8822_o;
  reg n8823_o;
  wire n8824_o;
  reg n8825_o;
  wire [31:0] n8827_o;
  wire n8828_o;
  wire n8829_o;
  wire [31:0] n8830_o;
  wire [31:0] n8831_o;
  wire n8832_o;
  wire n8833_o;
  wire n8834_o;
  wire n8835_o;
  wire n8836_o;
  wire n8837_o;
  wire n8838_o;
  wire n8839_o;
  wire n8840_o;
  wire n8841_o;
  wire n8842_o;
  wire n8843_o;
  wire n8844_o;
  wire n8845_o;
  wire n8846_o;
  wire n8847_o;
  wire n8848_o;
  wire n8849_o;
  wire n8850_o;
  wire n8851_o;
  wire n8852_o;
  wire n8853_o;
  wire n8854_o;
  wire [31:0] n8855_o;
  wire [31:0] n8857_o;
  wire [31:0] n8858_o;
  wire [31:0] n8860_o;
  wire [31:0] n8861_o;
  wire n8862_o;
  wire n8863_o;
  wire [31:0] n8864_o;
  wire [31:0] n8865_o;
  wire [3:0] n8866_o;
  wire [3:0] n8868_o;
  wire [3:0] n8869_o;
  wire [3:0] n8871_o;
  wire [3:0] n8872_o;
  wire n8873_o;
  wire n8874_o;
  wire [3:0] n8875_o;
  wire [3:0] n8876_o;
  wire n8877_o;
  wire [31:0] n8878_o;
  wire n8879_o;
  wire n8880_o;
  wire n8881_o;
  wire n8882_o;
  wire n8884_o;
  wire n8885_o;
  wire n8886_o;
  wire n8887_o;
  wire [31:0] n8889_o;
  wire n8890_o;
  wire n8891_o;
  wire n8892_o;
  wire n8894_o;
  wire n8895_o;
  wire n8896_o;
  reg [1:0] n8898_q;
  reg [1:0] n8899_q;
  wire [7:0] n8900_o;
  wire [33:0] n8901_o;
  wire [33:0] n8902_o;
  wire [73:0] n8903_o;
  assign a_rsp_o_data = n8735_o; //(module output)
  assign a_rsp_o_ack = n8736_o; //(module output)
  assign a_rsp_o_err = n8737_o; //(module output)
  assign b_rsp_o_data = n8740_o; //(module output)
  assign b_rsp_o_ack = n8741_o; //(module output)
  assign b_rsp_o_err = n8742_o; //(module output)
  assign x_req_o_addr = n8744_o; //(module output)
  assign x_req_o_data = n8745_o; //(module output)
  assign x_req_o_ben = n8746_o; //(module output)
  assign x_req_o_stb = n8747_o; //(module output)
  assign x_req_o_rw = n8748_o; //(module output)
  assign x_req_o_src = n8749_o; //(module output)
  assign x_req_o_priv = n8750_o; //(module output)
  assign x_req_o_rvso = n8751_o; //(module output)
  assign x_req_o_fence = n8752_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:875:5  */
  assign n8733_o = {a_req_i_fence, a_req_i_rvso, a_req_i_priv, a_req_i_src, a_req_i_rw, a_req_i_stb, a_req_i_ben, a_req_i_data, a_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:873:5  */
  assign n8735_o = n8901_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:872:5  */
  assign n8736_o = n8901_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:868:5  */
  assign n8737_o = n8901_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:867:5  */
  assign n8738_o = {b_req_i_fence, b_req_i_rvso, b_req_i_priv, b_req_i_src, b_req_i_rw, b_req_i_stb, b_req_i_ben, b_req_i_data, b_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:860:5  */
  assign n8740_o = n8902_o[31:0]; // extract
  assign n8741_o = n8902_o[32]; // extract
  assign n8742_o = n8902_o[33]; // extract
  assign n8744_o = n8903_o[31:0]; // extract
  assign n8745_o = n8903_o[63:32]; // extract
  assign n8746_o = n8903_o[67:64]; // extract
  assign n8747_o = n8903_o[68]; // extract
  assign n8748_o = n8903_o[69]; // extract
  assign n8749_o = n8903_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1034:14  */
  assign n8750_o = n8903_o[71]; // extract
  assign n8751_o = n8903_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:717:12  */
  assign n8752_o = n8903_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:717:12  */
  assign n8753_o = {x_rsp_i_err, x_rsp_i_ack, x_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:69:10  */
  assign arbiter = n8900_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:82:16  */
  assign n8755_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:87:32  */
  assign n8760_o = arbiter[3:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:33  */
  assign n8761_o = arbiter[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:50  */
  assign n8762_o = n8733_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:39  */
  assign n8763_o = n8761_o | n8762_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:77  */
  assign n8764_o = arbiter[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:60  */
  assign n8765_o = ~n8764_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:55  */
  assign n8766_o = n8763_o & n8765_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:33  */
  assign n8767_o = arbiter[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:50  */
  assign n8768_o = n8738_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:39  */
  assign n8769_o = n8767_o | n8768_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:77  */
  assign n8770_o = arbiter[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:60  */
  assign n8771_o = ~n8770_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:55  */
  assign n8772_o = n8769_o & n8771_o;
  assign n8773_o = {n8772_o, n8766_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:936:3  */
  assign n8778_o = {1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:97:34  */
  assign n8783_o = arbiter[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:102:18  */
  assign n8786_o = arbiter[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:107:21  */
  assign n8788_o = n8753_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:107:44  */
  assign n8789_o = n8753_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:107:32  */
  assign n8790_o = n8788_o | n8789_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:107:9  */
  assign n8791_o = n8790_o ? 2'b00 : n8783_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:104:7  */
  assign n8793_o = n8786_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:114:21  */
  assign n8795_o = n8753_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:114:44  */
  assign n8796_o = n8753_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:114:32  */
  assign n8797_o = n8795_o | n8796_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:114:9  */
  assign n8798_o = n8797_o ? 2'b00 : n8783_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:111:7  */
  assign n8800_o = n8786_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:21  */
  assign n8801_o = n8733_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:44  */
  assign n8802_o = arbiter[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:32  */
  assign n8803_o = n8801_o | n8802_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:24  */
  assign n8807_o = n8738_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:47  */
  assign n8808_o = arbiter[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:35  */
  assign n8809_o = n8807_o | n8808_o;
  assign n8813_o = {1'b1, 1'b1};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:9  */
  assign n8814_o = n8809_o ? 2'b10 : n8783_o;
  assign n8815_o = {1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:9  */
  assign n8816_o = n8809_o ? n8813_o : n8815_o;
  assign n8817_o = {1'b1, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:9  */
  assign n8818_o = n8803_o ? 2'b01 : n8814_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:9  */
  assign n8819_o = n8803_o ? n8817_o : n8816_o;
  assign n8820_o = {n8800_o, n8793_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:102:5  */
  always @*
    case (n8820_o)
      2'b10: n8821_o = n8798_o;
      2'b01: n8821_o = n8791_o;
      default: n8821_o = n8818_o;
    endcase
  assign n8822_o = n8819_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:102:5  */
  always @*
    case (n8820_o)
      2'b10: n8823_o = 1'b1;
      2'b01: n8823_o = 1'b0;
      default: n8823_o = n8822_o;
    endcase
  assign n8824_o = n8819_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:102:5  */
  always @*
    case (n8820_o)
      2'b10: n8825_o = 1'b0;
      2'b01: n8825_o = 1'b0;
      default: n8825_o = n8824_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:28  */
  assign n8827_o = n8733_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:47  */
  assign n8828_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:51  */
  assign n8829_o = ~n8828_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:33  */
  assign n8830_o = n8829_o ? n8827_o : n8831_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:71  */
  assign n8831_o = n8738_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:28  */
  assign n8832_o = n8733_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:47  */
  assign n8833_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:51  */
  assign n8834_o = ~n8833_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:33  */
  assign n8835_o = n8834_o ? n8832_o : n8836_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:71  */
  assign n8836_o = n8738_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:28  */
  assign n8837_o = n8733_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:47  */
  assign n8838_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:51  */
  assign n8839_o = ~n8838_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:33  */
  assign n8840_o = n8839_o ? n8837_o : n8841_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:71  */
  assign n8841_o = n8738_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:28  */
  assign n8842_o = n8733_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:47  */
  assign n8843_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:51  */
  assign n8844_o = ~n8843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:33  */
  assign n8845_o = n8844_o ? n8842_o : n8846_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:71  */
  assign n8846_o = n8738_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:28  */
  assign n8847_o = n8733_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:47  */
  assign n8848_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:51  */
  assign n8849_o = ~n8848_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:33  */
  assign n8850_o = n8849_o ? n8847_o : n8851_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:71  */
  assign n8851_o = n8738_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:141:28  */
  assign n8852_o = n8733_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:141:45  */
  assign n8853_o = n8738_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:141:34  */
  assign n8854_o = n8852_o | n8853_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:143:28  */
  assign n8855_o = n8738_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:143:33  */
  assign n8857_o = 1'b0 ? n8855_o : n8860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:144:28  */
  assign n8858_o = n8733_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:143:58  */
  assign n8860_o = 1'b0 ? n8858_o : n8864_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:145:28  */
  assign n8861_o = n8733_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:145:47  */
  assign n8862_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:145:51  */
  assign n8863_o = ~n8862_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:144:58  */
  assign n8864_o = n8863_o ? n8861_o : n8865_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:145:71  */
  assign n8865_o = n8738_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:147:28  */
  assign n8866_o = n8738_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:147:32  */
  assign n8868_o = 1'b0 ? n8866_o : n8871_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:148:28  */
  assign n8869_o = n8733_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:147:58  */
  assign n8871_o = 1'b0 ? n8869_o : n8875_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:149:28  */
  assign n8872_o = n8733_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:149:46  */
  assign n8873_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:149:50  */
  assign n8874_o = ~n8873_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:148:58  */
  assign n8875_o = n8874_o ? n8872_o : n8876_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:149:71  */
  assign n8876_o = n8738_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:151:28  */
  assign n8877_o = arbiter[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:156:27  */
  assign n8878_o = n8753_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:157:27  */
  assign n8879_o = n8753_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:157:45  */
  assign n8880_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:157:49  */
  assign n8881_o = ~n8880_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:157:31  */
  assign n8882_o = n8881_o ? n8879_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:158:27  */
  assign n8884_o = n8753_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:158:45  */
  assign n8885_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:158:49  */
  assign n8886_o = ~n8885_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:158:31  */
  assign n8887_o = n8886_o ? n8884_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:160:27  */
  assign n8889_o = n8753_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:161:27  */
  assign n8890_o = n8753_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:161:45  */
  assign n8891_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:161:31  */
  assign n8892_o = n8891_o ? n8890_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:162:27  */
  assign n8894_o = n8753_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:162:45  */
  assign n8895_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:162:31  */
  assign n8896_o = n8895_o ? n8894_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:86:5  */
  always @(posedge clk_i or posedge n8755_o)
    if (n8755_o)
      n8898_q <= n8778_o;
    else
      n8898_q <= n8773_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:86:5  */
  always @(posedge clk_i or posedge n8755_o)
    if (n8755_o)
      n8899_q <= 2'b00;
    else
      n8899_q <= n8760_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:82:5  */
  assign n8900_o = {n8825_o, n8823_o, n8898_q, n8821_o, n8899_q};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:82:5  */
  assign n8901_o = {n8887_o, n8882_o, n8878_o};
  assign n8902_o = {n8896_o, n8892_o, n8889_o};
  assign n8903_o = {n8854_o, n8835_o, n8840_o, n8845_o, n8850_o, n8877_o, n8868_o, n8857_o, n8830_o};
endmodule

module neorv32_cache_bus_32_32_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  rstn_i,
   input  clk_i,
   input  [31:0] host_req_i_addr,
   input  [31:0] host_req_i_data,
   input  [3:0] host_req_i_ben,
   input  host_req_i_stb,
   input  host_req_i_rw,
   input  host_req_i_src,
   input  host_req_i_priv,
   input  host_req_i_rvso,
   input  host_req_i_fence,
   input  [31:0] bus_rsp_i_data,
   input  bus_rsp_i_ack,
   input  bus_rsp_i_err,
   input  cmd_sync_i,
   input  cmd_miss_i,
   input  dirty_i,
   input  [31:0] base_i,
   input  [31:0] rdata_i,
   output [31:0] bus_req_o_addr,
   output [31:0] bus_req_o_data,
   output [3:0] bus_req_o_ben,
   output bus_req_o_stb,
   output bus_req_o_rw,
   output bus_req_o_src,
   output bus_req_o_priv,
   output bus_req_o_rvso,
   output bus_req_o_fence,
   output cmd_busy_o,
   output inval_o,
   output new_o,
   output [31:0] addr_o,
   output [3:0] we_o,
   output swe_o,
   output [31:0] wdata_o,
   output wstat_o);
  wire [73:0] n8472_o;
  wire [31:0] n8474_o;
  wire [31:0] n8475_o;
  wire [3:0] n8476_o;
  wire n8477_o;
  wire n8478_o;
  wire n8479_o;
  wire n8480_o;
  wire n8481_o;
  wire n8482_o;
  wire [33:0] n8483_o;
  wire [3:0] state;
  wire [3:0] upret;
  wire [3:0] state_nxt;
  wire [3:0] upret_nxt;
  wire [29:0] haddr;
  wire [29:0] baddr;
  wire [29:0] addr;
  wire [29:0] addr_nxt;
  wire [21:0] n8492_o;
  wire [21:0] n8495_o;
  wire [4:0] n8496_o;
  wire n8499_o;
  wire [29:0] n8511_o;
  wire [21:0] n8515_o;
  wire [4:0] n8516_o;
  wire [26:0] n8517_o;
  wire [2:0] n8518_o;
  wire [29:0] n8519_o;
  wire [31:0] n8521_o;
  wire [31:0] n8522_o;
  wire n8523_o;
  wire [21:0] n8524_o;
  wire [4:0] n8525_o;
  wire [26:0] n8526_o;
  wire [2:0] n8527_o;
  wire [29:0] n8528_o;
  wire [31:0] n8530_o;
  localparam [73:0] n8531_o = 74'b00000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [3:0] n8543_o;
  wire [3:0] n8545_o;
  wire n8547_o;
  wire [4:0] n8548_o;
  wire n8550_o;
  wire [21:0] n8551_o;
  wire [21:0] n8552_o;
  wire [3:0] n8555_o;
  wire [21:0] n8556_o;
  wire n8558_o;
  wire n8562_o;
  wire n8564_o;
  wire n8565_o;
  wire n8566_o;
  wire [2:0] n8567_o;
  wire [2:0] n8569_o;
  wire n8577_o;
  wire n8579_o;
  wire n8581_o;
  wire n8582_o;
  wire n8583_o;
  wire n8584_o;
  wire [3:0] n8587_o;
  wire [3:0] n8588_o;
  wire [2:0] n8589_o;
  wire [2:0] n8590_o;
  wire n8592_o;
  wire n8595_o;
  wire n8599_o;
  wire n8601_o;
  wire n8602_o;
  wire n8603_o;
  wire [2:0] n8604_o;
  wire [2:0] n8606_o;
  wire n8614_o;
  wire n8616_o;
  wire n8618_o;
  wire n8619_o;
  wire n8620_o;
  wire n8621_o;
  wire [3:0] n8623_o;
  wire [3:0] n8624_o;
  wire [2:0] n8625_o;
  wire [2:0] n8626_o;
  wire n8628_o;
  wire n8631_o;
  wire n8633_o;
  wire [21:0] n8634_o;
  wire n8636_o;
  wire [4:0] n8637_o;
  wire [4:0] n8639_o;
  wire n8647_o;
  wire n8649_o;
  wire n8651_o;
  wire n8652_o;
  wire n8653_o;
  wire n8654_o;
  wire n8655_o;
  wire n8656_o;
  wire n8657_o;
  wire n8658_o;
  wire n8660_o;
  wire n8661_o;
  wire [3:0] n8664_o;
  wire n8665_o;
  wire n8666_o;
  wire [3:0] n8668_o;
  wire [4:0] n8669_o;
  wire [4:0] n8670_o;
  wire n8672_o;
  wire [9:0] n8673_o;
  wire n8674_o;
  reg n8675_o;
  wire n8676_o;
  reg n8677_o;
  wire n8678_o;
  reg n8679_o;
  wire n8681_o;
  reg n8684_o;
  reg n8689_o;
  reg [3:0] n8693_o;
  reg n8697_o;
  reg [3:0] n8705_o;
  reg [3:0] n8708_o;
  wire [21:0] n8709_o;
  reg [21:0] n8710_o;
  wire [4:0] n8711_o;
  reg [4:0] n8712_o;
  wire [2:0] n8713_o;
  reg [2:0] n8714_o;
  wire n8720_o;
  wire n8722_o;
  wire n8723_o;
  wire n8724_o;
  reg [3:0] n8726_q;
  reg [3:0] n8727_q;
  wire [29:0] n8728_o;
  wire [29:0] n8729_o;
  reg [29:0] n8730_q;
  wire [29:0] n8731_o;
  wire [73:0] n8732_o;
  assign bus_req_o_addr = n8474_o; //(module output)
  assign bus_req_o_data = n8475_o; //(module output)
  assign bus_req_o_ben = n8476_o; //(module output)
  assign bus_req_o_stb = n8477_o; //(module output)
  assign bus_req_o_rw = n8478_o; //(module output)
  assign bus_req_o_src = n8479_o; //(module output)
  assign bus_req_o_priv = n8480_o; //(module output)
  assign bus_req_o_rvso = n8481_o; //(module output)
  assign bus_req_o_fence = n8482_o; //(module output)
  assign cmd_busy_o = n8724_o; //(module output)
  assign inval_o = n8684_o; //(module output)
  assign new_o = n8689_o; //(module output)
  assign addr_o = n8521_o; //(module output)
  assign we_o = n8693_o; //(module output)
  assign swe_o = n8697_o; //(module output)
  assign wdata_o = n8522_o; //(module output)
  assign wstat_o = n8523_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:33  */
  assign n8472_o = {host_req_i_fence, host_req_i_rvso, host_req_i_priv, host_req_i_src, host_req_i_rw, host_req_i_stb, host_req_i_ben, host_req_i_data, host_req_i_addr};
  assign n8474_o = n8732_o[31:0]; // extract
  assign n8475_o = n8732_o[63:32]; // extract
  assign n8476_o = n8732_o[67:64]; // extract
  assign n8477_o = n8732_o[68]; // extract
  assign n8478_o = n8732_o[69]; // extract
  assign n8479_o = n8732_o[70]; // extract
  assign n8480_o = n8732_o[71]; // extract
  assign n8481_o = n8732_o[72]; // extract
  assign n8482_o = n8732_o[73]; // extract
  assign n8483_o = {bus_rsp_i_err, bus_rsp_i_ack, bus_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:891:10  */
  assign state = n8726_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:891:17  */
  assign upret = n8727_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:891:24  */
  assign state_nxt = n8705_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:891:35  */
  assign upret_nxt = n8708_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:899:10  */
  assign haddr = n8728_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:899:17  */
  assign baddr = n8729_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:899:24  */
  assign addr = n8730_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:899:30  */
  assign addr_nxt = n8731_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:906:31  */
  assign n8492_o = n8472_o[31:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:911:22  */
  assign n8495_o = base_i[31:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:912:22  */
  assign n8496_o = base_i[9:5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:920:16  */
  assign n8499_o = ~rstn_i;
  assign n8511_o = {3'b000, 5'b00000, 22'b0000000000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:944:21  */
  assign n8515_o = addr[21:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:944:32  */
  assign n8516_o = addr[26:22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:944:25  */
  assign n8517_o = {n8515_o, n8516_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:944:43  */
  assign n8518_o = addr[29:27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:944:36  */
  assign n8519_o = {n8517_o, n8518_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:944:47  */
  assign n8521_o = {n8519_o, 2'b00};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:947:26  */
  assign n8522_o = n8483_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:948:26  */
  assign n8523_o = n8483_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:956:28  */
  assign n8524_o = addr[21:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:956:39  */
  assign n8525_o = addr[26:22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:956:32  */
  assign n8526_o = {n8524_o, n8525_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:956:50  */
  assign n8527_o = addr[29:27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:956:43  */
  assign n8528_o = {n8526_o, n8527_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:956:54  */
  assign n8530_o = {n8528_o, 2'b00};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:970:9  */
  assign n8543_o = cmd_miss_i ? 4'b0001 : state;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:968:9  */
  assign n8545_o = cmd_sync_i ? 4'b0111 : n8543_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:965:7  */
  assign n8547_o = state == 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:977:31  */
  assign n8548_o = baddr[26:22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:978:28  */
  assign n8550_o = 1'b1 & dirty_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:979:33  */
  assign n8551_o = baddr[21:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:982:33  */
  assign n8552_o = haddr[21:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:978:9  */
  assign n8555_o = n8550_o ? 4'b0100 : 4'b0010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:978:9  */
  assign n8556_o = n8550_o ? n8551_o : n8552_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:974:7  */
  assign n8558_o = state == 4'b0001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:987:7  */
  assign n8562_o = state == 4'b0010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:999:23  */
  assign n8564_o = n8483_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:999:48  */
  assign n8565_o = n8483_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:999:34  */
  assign n8566_o = n8564_o | n8565_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1000:59  */
  assign n8567_o = addr[29:27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1000:64  */
  assign n8569_o = n8567_o + 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8577_o = addr[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8579_o = 1'b1 & n8577_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8581_o = addr[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8582_o = n8579_o & n8581_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8583_o = addr[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8584_o = n8582_o & n8583_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1001:11  */
  assign n8587_o = n8584_o ? 4'b0000 : 4'b0010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:999:9  */
  assign n8588_o = n8566_o ? n8587_o : state;
  assign n8589_o = addr[29:27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:999:9  */
  assign n8590_o = n8566_o ? n8569_o : n8589_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:993:7  */
  assign n8592_o = state == 4'b0011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1009:7  */
  assign n8595_o = state == 4'b0100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1018:7  */
  assign n8599_o = state == 4'b0101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1035:25  */
  assign n8601_o = n8483_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1035:50  */
  assign n8602_o = n8483_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1035:36  */
  assign n8603_o = n8601_o | n8602_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1036:61  */
  assign n8604_o = addr[29:27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1036:66  */
  assign n8606_o = n8604_o + 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8614_o = addr[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8616_o = 1'b1 & n8614_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8618_o = addr[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8619_o = n8616_o & n8618_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8620_o = addr[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8621_o = n8619_o & n8620_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1037:13  */
  assign n8623_o = n8621_o ? upret : 4'b0100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1035:11  */
  assign n8624_o = n8603_o ? n8623_o : state;
  assign n8625_o = addr[29:27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1035:11  */
  assign n8626_o = n8603_o ? n8606_o : n8625_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1028:7  */
  assign n8628_o = state == 4'b0110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1046:7  */
  assign n8631_o = state == 4'b0111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1052:7  */
  assign n8633_o = state == 4'b1000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1058:31  */
  assign n8634_o = baddr[21:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1060:28  */
  assign n8636_o = 1'b1 & dirty_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1063:59  */
  assign n8637_o = addr[26:22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1063:64  */
  assign n8639_o = n8637_o + 5'b00001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8647_o = addr[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8649_o = 1'b1 & n8647_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8651_o = addr[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8652_o = n8649_o & n8651_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8653_o = addr[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8654_o = n8652_o & n8653_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8655_o = addr[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8656_o = n8654_o & n8655_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n8657_o = addr[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n8658_o = n8656_o & n8657_o;
  assign n8660_o = n8531_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1064:11  */
  assign n8661_o = n8658_o ? 1'b1 : n8660_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1064:11  */
  assign n8664_o = n8658_o ? 4'b0000 : 4'b1000;
  assign n8665_o = n8531_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1060:9  */
  assign n8666_o = n8636_o ? n8665_o : n8661_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1060:9  */
  assign n8668_o = n8636_o ? 4'b0100 : n8664_o;
  assign n8669_o = addr[26:22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1060:9  */
  assign n8670_o = n8636_o ? n8669_o : n8639_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1056:7  */
  assign n8672_o = state == 4'b1001;
  assign n8673_o = {n8672_o, n8633_o, n8631_o, n8628_o, n8599_o, n8595_o, n8592_o, n8562_o, n8558_o, n8547_o};
  assign n8674_o = n8531_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8675_o = n8674_o;
      10'b0100000000: n8675_o = n8674_o;
      10'b0010000000: n8675_o = n8674_o;
      10'b0001000000: n8675_o = n8674_o;
      10'b0000100000: n8675_o = 1'b1;
      10'b0000010000: n8675_o = n8674_o;
      10'b0000001000: n8675_o = n8674_o;
      10'b0000000100: n8675_o = 1'b1;
      10'b0000000010: n8675_o = n8674_o;
      10'b0000000001: n8675_o = n8674_o;
      default: n8675_o = n8674_o;
    endcase
  assign n8676_o = n8531_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8677_o = n8676_o;
      10'b0100000000: n8677_o = n8676_o;
      10'b0010000000: n8677_o = n8676_o;
      10'b0001000000: n8677_o = 1'b1;
      10'b0000100000: n8677_o = 1'b1;
      10'b0000010000: n8677_o = 1'b1;
      10'b0000001000: n8677_o = 1'b0;
      10'b0000000100: n8677_o = 1'b0;
      10'b0000000010: n8677_o = n8676_o;
      10'b0000000001: n8677_o = n8676_o;
      default: n8677_o = n8676_o;
    endcase
  assign n8678_o = n8531_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8679_o = n8666_o;
      10'b0100000000: n8679_o = n8678_o;
      10'b0010000000: n8679_o = n8678_o;
      10'b0001000000: n8679_o = n8678_o;
      10'b0000100000: n8679_o = n8678_o;
      10'b0000010000: n8679_o = n8678_o;
      10'b0000001000: n8679_o = n8678_o;
      10'b0000000100: n8679_o = n8678_o;
      10'b0000000010: n8679_o = n8678_o;
      10'b0000000001: n8679_o = n8678_o;
      default: n8679_o = n8678_o;
    endcase
  assign n8681_o = n8531_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8684_o = 1'b1;
      10'b0100000000: n8684_o = 1'b0;
      10'b0010000000: n8684_o = 1'b0;
      10'b0001000000: n8684_o = 1'b0;
      10'b0000100000: n8684_o = 1'b0;
      10'b0000010000: n8684_o = 1'b0;
      10'b0000001000: n8684_o = 1'b0;
      10'b0000000100: n8684_o = 1'b0;
      10'b0000000010: n8684_o = 1'b0;
      10'b0000000001: n8684_o = 1'b0;
      default: n8684_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8689_o = 1'b0;
      10'b0100000000: n8689_o = 1'b0;
      10'b0010000000: n8689_o = 1'b0;
      10'b0001000000: n8689_o = 1'b1;
      10'b0000100000: n8689_o = 1'b0;
      10'b0000010000: n8689_o = 1'b0;
      10'b0000001000: n8689_o = 1'b1;
      10'b0000000100: n8689_o = 1'b0;
      10'b0000000010: n8689_o = 1'b0;
      10'b0000000001: n8689_o = 1'b0;
      default: n8689_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8693_o = 4'b0000;
      10'b0100000000: n8693_o = 4'b0000;
      10'b0010000000: n8693_o = 4'b0000;
      10'b0001000000: n8693_o = 4'b0000;
      10'b0000100000: n8693_o = 4'b0000;
      10'b0000010000: n8693_o = 4'b0000;
      10'b0000001000: n8693_o = 4'b1111;
      10'b0000000100: n8693_o = 4'b0000;
      10'b0000000010: n8693_o = 4'b0000;
      10'b0000000001: n8693_o = 4'b0000;
      default: n8693_o = 4'b0000;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8697_o = 1'b0;
      10'b0100000000: n8697_o = 1'b0;
      10'b0010000000: n8697_o = 1'b0;
      10'b0001000000: n8697_o = 1'b0;
      10'b0000100000: n8697_o = 1'b0;
      10'b0000010000: n8697_o = 1'b0;
      10'b0000001000: n8697_o = 1'b1;
      10'b0000000100: n8697_o = 1'b0;
      10'b0000000010: n8697_o = 1'b0;
      10'b0000000001: n8697_o = 1'b0;
      default: n8697_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8705_o = n8668_o;
      10'b0100000000: n8705_o = 4'b1001;
      10'b0010000000: n8705_o = 4'b1000;
      10'b0001000000: n8705_o = n8624_o;
      10'b0000100000: n8705_o = 4'b0110;
      10'b0000010000: n8705_o = 4'b0101;
      10'b0000001000: n8705_o = n8588_o;
      10'b0000000100: n8705_o = 4'b0011;
      10'b0000000010: n8705_o = n8555_o;
      10'b0000000001: n8705_o = n8545_o;
      default: n8705_o = 4'b0000;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8708_o = upret;
      10'b0100000000: n8708_o = upret;
      10'b0010000000: n8708_o = 4'b1001;
      10'b0001000000: n8708_o = upret;
      10'b0000100000: n8708_o = upret;
      10'b0000010000: n8708_o = upret;
      10'b0000001000: n8708_o = upret;
      10'b0000000100: n8708_o = upret;
      10'b0000000010: n8708_o = 4'b0010;
      10'b0000000001: n8708_o = upret;
      default: n8708_o = upret;
    endcase
  assign n8709_o = addr[21:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8710_o = n8634_o;
      10'b0100000000: n8710_o = n8709_o;
      10'b0010000000: n8710_o = n8709_o;
      10'b0001000000: n8710_o = n8709_o;
      10'b0000100000: n8710_o = n8709_o;
      10'b0000010000: n8710_o = n8709_o;
      10'b0000001000: n8710_o = n8709_o;
      10'b0000000100: n8710_o = n8709_o;
      10'b0000000010: n8710_o = n8556_o;
      10'b0000000001: n8710_o = n8709_o;
      default: n8710_o = n8709_o;
    endcase
  assign n8711_o = addr[26:22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8712_o = n8670_o;
      10'b0100000000: n8712_o = n8711_o;
      10'b0010000000: n8712_o = 5'b00000;
      10'b0001000000: n8712_o = n8711_o;
      10'b0000100000: n8712_o = n8711_o;
      10'b0000010000: n8712_o = n8711_o;
      10'b0000001000: n8712_o = n8711_o;
      10'b0000000100: n8712_o = n8711_o;
      10'b0000000010: n8712_o = n8548_o;
      10'b0000000001: n8712_o = n8711_o;
      default: n8712_o = n8711_o;
    endcase
  assign n8713_o = addr[29:27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:963:5  */
  always @*
    case (n8673_o)
      10'b1000000000: n8714_o = n8713_o;
      10'b0100000000: n8714_o = n8713_o;
      10'b0010000000: n8714_o = n8713_o;
      10'b0001000000: n8714_o = n8626_o;
      10'b0000100000: n8714_o = n8713_o;
      10'b0000010000: n8714_o = n8713_o;
      10'b0000001000: n8714_o = n8590_o;
      10'b0000000100: n8714_o = n8713_o;
      10'b0000000010: n8714_o = n8713_o;
      10'b0000000001: n8714_o = 3'b000;
      default: n8714_o = n8713_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1081:33  */
  assign n8720_o = state == 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1081:53  */
  assign n8722_o = state == 4'b0001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1081:43  */
  assign n8723_o = n8720_o | n8722_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:1081:21  */
  assign n8724_o = n8723_o ? 1'b0 : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:926:5  */
  always @(posedge clk_i or posedge n8499_o)
    if (n8499_o)
      n8726_q <= 4'b0000;
    else
      n8726_q <= state_nxt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:926:5  */
  always @(posedge clk_i or posedge n8499_o)
    if (n8499_o)
      n8727_q <= 4'b0000;
    else
      n8727_q <= upret_nxt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:920:5  */
  assign n8728_o = {3'b000, 5'b00000, n8492_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:920:5  */
  assign n8729_o = {3'b000, n8496_o, n8495_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:926:5  */
  always @(posedge clk_i or posedge n8499_o)
    if (n8499_o)
      n8730_q <= n8511_o;
    else
      n8730_q <= addr_nxt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:920:5  */
  assign n8731_o = {n8714_o, n8712_o, n8710_o};
  assign n8732_o = {n8679_o, n8681_o, 1'b0, 1'b0, n8677_o, n8675_o, 4'b1111, rdata_i, n8530_o};
endmodule

module neorv32_cache_memory_32_32_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  rstn_i,
   input  clk_i,
   input  inval_i,
   input  new_i,
   input  dirty_i,
   input  [31:0] addr_i,
   input  [3:0] we_i,
   input  swe_i,
   input  [31:0] wdata_i,
   input  wstat_i,
   output hit_o,
   output dirty_o,
   output [31:0] base_o,
   output [31:0] rdata_o,
   output rstat_o);
  wire [31:0] valid_mem;
  wire [31:0] dirty_mem;
  wire valid_mem_rd;
  wire dirty_mem_rd;
  wire [21:0] tag_mem_rd;
  wire [31:0] data_mem_rd;
  wire stat_mem_rd;
  wire [21:0] acc_tag;
  wire [21:0] acc_tag_ff;
  wire [4:0] acc_idx;
  wire [4:0] acc_idx_ff;
  wire [2:0] acc_off;
  wire [7:0] acc_adr;
  wire [21:0] n7623_o;
  wire [4:0] n7624_o;
  wire [2:0] n7625_o;
  wire [7:0] n7626_o;
  wire n7628_o;
  wire n7638_o;
  wire [31:0] n7652_o;
  wire [31:0] n7657_o;
  wire [31:0] n7658_o;
  wire [31:0] n7659_o;
  wire n7694_o;
  wire n7695_o;
  wire n7696_o;
  wire n7699_o;
  wire n7701_o;
  wire n7702_o;
  wire n7707_o;
  wire [7:0] n7712_o;
  wire n7715_o;
  wire [7:0] n7720_o;
  wire n7723_o;
  wire [7:0] n7728_o;
  wire n7731_o;
  wire [7:0] n7736_o;
  wire [31:0] n7770_o;
  wire n7775_o;
  reg [31:0] n7776_q;
  reg [31:0] n7777_q;
  wire n7778_o;
  wire n7779_o;
  reg n7780_q;
  wire n7781_o;
  wire n7782_o;
  reg n7783_q;
  reg [21:0] n7799_q;
  reg [4:0] n7800_q;
  wire [31:0] n7801_o;
  reg [21:0] n7803_data; // mem_rd
  reg [7:0] n7810_data; // mem_rd
  reg [7:0] n7813_data; // mem_rd
  reg [7:0] n7816_data; // mem_rd
  reg [7:0] n7819_data; // mem_rd
  reg n7822_data; // mem_rd
  wire n7824_o;
  wire n7825_o;
  wire n7826_o;
  wire n7827_o;
  wire n7828_o;
  wire n7829_o;
  wire n7830_o;
  wire n7831_o;
  wire n7832_o;
  wire n7833_o;
  wire n7834_o;
  wire n7835_o;
  wire n7836_o;
  wire n7837_o;
  wire n7838_o;
  wire n7839_o;
  wire n7840_o;
  wire n7841_o;
  wire n7842_o;
  wire n7843_o;
  wire n7844_o;
  wire n7845_o;
  wire n7846_o;
  wire n7847_o;
  wire n7848_o;
  wire n7849_o;
  wire n7850_o;
  wire n7851_o;
  wire n7852_o;
  wire n7853_o;
  wire n7854_o;
  wire n7855_o;
  wire n7856_o;
  wire n7857_o;
  wire n7858_o;
  wire n7859_o;
  wire n7860_o;
  wire n7861_o;
  wire n7862_o;
  wire n7863_o;
  wire n7864_o;
  wire n7865_o;
  wire n7866_o;
  wire n7867_o;
  wire n7868_o;
  wire n7869_o;
  wire n7870_o;
  wire n7871_o;
  wire n7872_o;
  wire n7873_o;
  wire n7874_o;
  wire n7875_o;
  wire n7876_o;
  wire n7877_o;
  wire n7878_o;
  wire n7879_o;
  wire n7880_o;
  wire n7881_o;
  wire n7882_o;
  wire n7883_o;
  wire n7884_o;
  wire n7885_o;
  wire n7886_o;
  wire n7887_o;
  wire n7888_o;
  wire n7889_o;
  wire n7890_o;
  wire n7891_o;
  wire n7892_o;
  wire n7893_o;
  wire n7894_o;
  wire n7895_o;
  wire n7896_o;
  wire n7897_o;
  wire n7898_o;
  wire n7899_o;
  wire n7900_o;
  wire n7901_o;
  wire n7902_o;
  wire n7903_o;
  wire n7904_o;
  wire n7905_o;
  wire n7906_o;
  wire n7907_o;
  wire n7908_o;
  wire n7909_o;
  wire n7910_o;
  wire n7911_o;
  wire n7912_o;
  wire n7913_o;
  wire n7914_o;
  wire n7915_o;
  wire n7916_o;
  wire n7917_o;
  wire n7918_o;
  wire n7919_o;
  wire n7920_o;
  wire n7921_o;
  wire n7922_o;
  wire n7923_o;
  wire n7924_o;
  wire n7925_o;
  wire n7926_o;
  wire n7927_o;
  wire n7928_o;
  wire n7929_o;
  wire n7930_o;
  wire n7931_o;
  wire n7932_o;
  wire n7933_o;
  wire n7934_o;
  wire n7935_o;
  wire n7936_o;
  wire n7937_o;
  wire n7938_o;
  wire n7939_o;
  wire n7940_o;
  wire n7941_o;
  wire n7942_o;
  wire n7943_o;
  wire n7944_o;
  wire n7945_o;
  wire n7946_o;
  wire n7947_o;
  wire n7948_o;
  wire n7949_o;
  wire n7950_o;
  wire n7951_o;
  wire n7952_o;
  wire n7953_o;
  wire n7954_o;
  wire n7955_o;
  wire n7956_o;
  wire n7957_o;
  wire [31:0] n7958_o;
  wire n7959_o;
  wire n7960_o;
  wire n7961_o;
  wire n7962_o;
  wire n7963_o;
  wire n7964_o;
  wire n7965_o;
  wire n7966_o;
  wire n7967_o;
  wire n7968_o;
  wire n7969_o;
  wire n7970_o;
  wire n7971_o;
  wire n7972_o;
  wire n7973_o;
  wire n7974_o;
  wire n7975_o;
  wire n7976_o;
  wire n7977_o;
  wire n7978_o;
  wire n7979_o;
  wire n7980_o;
  wire n7981_o;
  wire n7982_o;
  wire n7983_o;
  wire n7984_o;
  wire n7985_o;
  wire n7986_o;
  wire n7987_o;
  wire n7988_o;
  wire n7989_o;
  wire n7990_o;
  wire n7991_o;
  wire n7992_o;
  wire n7993_o;
  wire n7994_o;
  wire n7995_o;
  wire n7996_o;
  wire n7997_o;
  wire n7998_o;
  wire n7999_o;
  wire n8000_o;
  wire n8001_o;
  wire n8002_o;
  wire n8003_o;
  wire n8004_o;
  wire n8005_o;
  wire n8006_o;
  wire n8007_o;
  wire n8008_o;
  wire n8009_o;
  wire n8010_o;
  wire n8011_o;
  wire n8012_o;
  wire n8013_o;
  wire n8014_o;
  wire n8015_o;
  wire n8016_o;
  wire n8017_o;
  wire n8018_o;
  wire n8019_o;
  wire n8020_o;
  wire n8021_o;
  wire n8022_o;
  wire n8023_o;
  wire n8024_o;
  wire n8025_o;
  wire n8026_o;
  wire n8027_o;
  wire n8028_o;
  wire n8029_o;
  wire n8030_o;
  wire n8031_o;
  wire n8032_o;
  wire n8033_o;
  wire n8034_o;
  wire n8035_o;
  wire n8036_o;
  wire n8037_o;
  wire n8038_o;
  wire n8039_o;
  wire n8040_o;
  wire n8041_o;
  wire n8042_o;
  wire n8043_o;
  wire n8044_o;
  wire n8045_o;
  wire n8046_o;
  wire n8047_o;
  wire n8048_o;
  wire n8049_o;
  wire n8050_o;
  wire n8051_o;
  wire n8052_o;
  wire n8053_o;
  wire n8054_o;
  wire n8055_o;
  wire n8056_o;
  wire n8057_o;
  wire n8058_o;
  wire n8059_o;
  wire n8060_o;
  wire n8061_o;
  wire n8062_o;
  wire n8063_o;
  wire n8064_o;
  wire n8065_o;
  wire n8066_o;
  wire n8067_o;
  wire n8068_o;
  wire n8069_o;
  wire n8070_o;
  wire n8071_o;
  wire n8072_o;
  wire n8073_o;
  wire n8074_o;
  wire n8075_o;
  wire n8076_o;
  wire n8077_o;
  wire n8078_o;
  wire n8079_o;
  wire n8080_o;
  wire n8081_o;
  wire n8082_o;
  wire n8083_o;
  wire n8084_o;
  wire n8085_o;
  wire n8086_o;
  wire n8087_o;
  wire n8088_o;
  wire n8089_o;
  wire n8090_o;
  wire n8091_o;
  wire n8092_o;
  wire [31:0] n8093_o;
  wire n8094_o;
  wire n8095_o;
  wire n8096_o;
  wire n8097_o;
  wire n8098_o;
  wire n8099_o;
  wire n8100_o;
  wire n8101_o;
  wire n8102_o;
  wire n8103_o;
  wire n8104_o;
  wire n8105_o;
  wire n8106_o;
  wire n8107_o;
  wire n8108_o;
  wire n8109_o;
  wire n8110_o;
  wire n8111_o;
  wire n8112_o;
  wire n8113_o;
  wire n8114_o;
  wire n8115_o;
  wire n8116_o;
  wire n8117_o;
  wire n8118_o;
  wire n8119_o;
  wire n8120_o;
  wire n8121_o;
  wire n8122_o;
  wire n8123_o;
  wire n8124_o;
  wire n8125_o;
  wire n8126_o;
  wire n8127_o;
  wire n8128_o;
  wire n8129_o;
  wire n8130_o;
  wire n8131_o;
  wire n8132_o;
  wire n8133_o;
  wire n8134_o;
  wire n8135_o;
  wire n8136_o;
  wire n8137_o;
  wire n8138_o;
  wire n8139_o;
  wire n8140_o;
  wire n8141_o;
  wire n8142_o;
  wire n8143_o;
  wire n8144_o;
  wire n8145_o;
  wire n8146_o;
  wire n8147_o;
  wire n8148_o;
  wire n8149_o;
  wire n8150_o;
  wire n8151_o;
  wire n8152_o;
  wire n8153_o;
  wire n8154_o;
  wire n8155_o;
  wire n8156_o;
  wire n8157_o;
  wire n8158_o;
  wire n8159_o;
  wire n8160_o;
  wire n8161_o;
  wire n8162_o;
  wire n8163_o;
  wire n8164_o;
  wire n8165_o;
  wire n8166_o;
  wire n8167_o;
  wire n8168_o;
  wire n8169_o;
  wire n8170_o;
  wire n8171_o;
  wire n8172_o;
  wire n8173_o;
  wire n8174_o;
  wire n8175_o;
  wire n8176_o;
  wire n8177_o;
  wire n8178_o;
  wire n8179_o;
  wire n8180_o;
  wire n8181_o;
  wire n8182_o;
  wire n8183_o;
  wire n8184_o;
  wire n8185_o;
  wire n8186_o;
  wire n8187_o;
  wire n8188_o;
  wire n8189_o;
  wire n8190_o;
  wire n8191_o;
  wire n8192_o;
  wire n8193_o;
  wire n8194_o;
  wire n8195_o;
  wire n8196_o;
  wire n8197_o;
  wire n8198_o;
  wire n8199_o;
  wire n8200_o;
  wire n8201_o;
  wire n8202_o;
  wire n8203_o;
  wire n8204_o;
  wire n8205_o;
  wire n8206_o;
  wire n8207_o;
  wire n8208_o;
  wire n8209_o;
  wire n8210_o;
  wire n8211_o;
  wire n8212_o;
  wire n8213_o;
  wire n8214_o;
  wire n8215_o;
  wire n8216_o;
  wire n8217_o;
  wire n8218_o;
  wire n8219_o;
  wire n8220_o;
  wire n8221_o;
  wire n8222_o;
  wire n8223_o;
  wire n8224_o;
  wire n8225_o;
  wire n8226_o;
  wire n8227_o;
  wire [31:0] n8228_o;
  wire n8229_o;
  wire n8230_o;
  wire n8231_o;
  wire n8232_o;
  wire n8233_o;
  wire n8234_o;
  wire n8235_o;
  wire n8236_o;
  wire n8237_o;
  wire n8238_o;
  wire n8239_o;
  wire n8240_o;
  wire n8241_o;
  wire n8242_o;
  wire n8243_o;
  wire n8244_o;
  wire n8245_o;
  wire n8246_o;
  wire n8247_o;
  wire n8248_o;
  wire n8249_o;
  wire n8250_o;
  wire n8251_o;
  wire n8252_o;
  wire n8253_o;
  wire n8254_o;
  wire n8255_o;
  wire n8256_o;
  wire n8257_o;
  wire n8258_o;
  wire n8259_o;
  wire n8260_o;
  wire n8261_o;
  wire n8262_o;
  wire n8263_o;
  wire n8264_o;
  wire n8265_o;
  wire n8266_o;
  wire n8267_o;
  wire n8268_o;
  wire n8269_o;
  wire n8270_o;
  wire n8271_o;
  wire n8272_o;
  wire n8273_o;
  wire n8274_o;
  wire n8275_o;
  wire n8276_o;
  wire n8277_o;
  wire n8278_o;
  wire n8279_o;
  wire n8280_o;
  wire n8281_o;
  wire n8282_o;
  wire n8283_o;
  wire n8284_o;
  wire n8285_o;
  wire n8286_o;
  wire n8287_o;
  wire n8288_o;
  wire n8289_o;
  wire n8290_o;
  wire n8291_o;
  wire n8292_o;
  wire n8293_o;
  wire n8294_o;
  wire n8295_o;
  wire n8296_o;
  wire n8297_o;
  wire n8298_o;
  wire n8299_o;
  wire n8300_o;
  wire n8301_o;
  wire n8302_o;
  wire n8303_o;
  wire n8304_o;
  wire n8305_o;
  wire n8306_o;
  wire n8307_o;
  wire n8308_o;
  wire n8309_o;
  wire n8310_o;
  wire n8311_o;
  wire n8312_o;
  wire n8313_o;
  wire n8314_o;
  wire n8315_o;
  wire n8316_o;
  wire n8317_o;
  wire n8318_o;
  wire n8319_o;
  wire n8320_o;
  wire n8321_o;
  wire n8322_o;
  wire n8323_o;
  wire n8324_o;
  wire n8325_o;
  wire n8326_o;
  wire n8327_o;
  wire n8328_o;
  wire n8329_o;
  wire n8330_o;
  wire n8331_o;
  wire n8332_o;
  wire n8333_o;
  wire n8334_o;
  wire n8335_o;
  wire n8336_o;
  wire n8337_o;
  wire n8338_o;
  wire n8339_o;
  wire n8340_o;
  wire n8341_o;
  wire n8342_o;
  wire n8343_o;
  wire n8344_o;
  wire n8345_o;
  wire n8346_o;
  wire n8347_o;
  wire n8348_o;
  wire n8349_o;
  wire n8350_o;
  wire n8351_o;
  wire n8352_o;
  wire n8353_o;
  wire n8354_o;
  wire n8355_o;
  wire n8356_o;
  wire n8357_o;
  wire n8358_o;
  wire n8359_o;
  wire n8360_o;
  wire n8361_o;
  wire n8362_o;
  wire [31:0] n8363_o;
  wire n8364_o;
  wire n8365_o;
  wire n8366_o;
  wire n8367_o;
  wire n8368_o;
  wire n8369_o;
  wire n8370_o;
  wire n8371_o;
  wire n8372_o;
  wire n8373_o;
  wire n8374_o;
  wire n8375_o;
  wire n8376_o;
  wire n8377_o;
  wire n8378_o;
  wire n8379_o;
  wire n8380_o;
  wire n8381_o;
  wire n8382_o;
  wire n8383_o;
  wire n8384_o;
  wire n8385_o;
  wire n8386_o;
  wire n8387_o;
  wire n8388_o;
  wire n8389_o;
  wire n8390_o;
  wire n8391_o;
  wire n8392_o;
  wire n8393_o;
  wire n8394_o;
  wire n8395_o;
  wire [1:0] n8396_o;
  reg n8397_o;
  wire [1:0] n8398_o;
  reg n8399_o;
  wire [1:0] n8400_o;
  reg n8401_o;
  wire [1:0] n8402_o;
  reg n8403_o;
  wire [1:0] n8404_o;
  reg n8405_o;
  wire [1:0] n8406_o;
  reg n8407_o;
  wire [1:0] n8408_o;
  reg n8409_o;
  wire [1:0] n8410_o;
  reg n8411_o;
  wire [1:0] n8412_o;
  reg n8413_o;
  wire [1:0] n8414_o;
  reg n8415_o;
  wire n8416_o;
  wire n8417_o;
  wire n8418_o;
  wire n8419_o;
  wire n8420_o;
  wire n8421_o;
  wire n8422_o;
  wire n8423_o;
  wire n8424_o;
  wire n8425_o;
  wire n8426_o;
  wire n8427_o;
  wire n8428_o;
  wire n8429_o;
  wire n8430_o;
  wire n8431_o;
  wire n8432_o;
  wire n8433_o;
  wire n8434_o;
  wire n8435_o;
  wire n8436_o;
  wire n8437_o;
  wire n8438_o;
  wire n8439_o;
  wire n8440_o;
  wire n8441_o;
  wire n8442_o;
  wire n8443_o;
  wire n8444_o;
  wire n8445_o;
  wire n8446_o;
  wire n8447_o;
  wire n8448_o;
  wire n8449_o;
  wire [1:0] n8450_o;
  reg n8451_o;
  wire [1:0] n8452_o;
  reg n8453_o;
  wire [1:0] n8454_o;
  reg n8455_o;
  wire [1:0] n8456_o;
  reg n8457_o;
  wire [1:0] n8458_o;
  reg n8459_o;
  wire [1:0] n8460_o;
  reg n8461_o;
  wire [1:0] n8462_o;
  reg n8463_o;
  wire [1:0] n8464_o;
  reg n8465_o;
  wire [1:0] n8466_o;
  reg n8467_o;
  wire [1:0] n8468_o;
  reg n8469_o;
  wire n8470_o;
  wire n8471_o;
  assign hit_o = n7696_o; //(module output)
  assign dirty_o = n7702_o; //(module output)
  assign base_o = n7801_o; //(module output)
  assign rdata_o = data_mem_rd; //(module output)
  assign rstat_o = n7775_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:670:10  */
  assign valid_mem = n7776_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:670:24  */
  assign dirty_mem = n7777_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:671:10  */
  assign valid_mem_rd = n7780_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:671:24  */
  assign dirty_mem_rd = n7783_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:676:10  */
  assign tag_mem_rd = n7803_data; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:681:10  */
  assign data_mem_rd = n7770_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:685:10  */
  assign stat_mem_rd = n7822_data; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:688:10  */
  assign acc_tag = n7623_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:688:19  */
  assign acc_tag_ff = n7799_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:689:10  */
  assign acc_idx = n7624_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:689:19  */
  assign acc_idx_ff = n7800_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:690:10  */
  assign acc_off = n7625_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:691:10  */
  assign acc_adr = n7626_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:697:20  */
  assign n7623_o = addr_i[31:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:698:20  */
  assign n7624_o = addr_i[9:5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:699:20  */
  assign n7625_o = addr_i[4:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:700:22  */
  assign n7626_o = {acc_idx, acc_off};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:705:16  */
  assign n7628_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:719:16  */
  assign n7638_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:727:9  */
  assign n7652_o = inval_i ? n8228_o : valid_mem;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:730:9  */
  assign n7657_o = dirty_i ? n8363_o : dirty_mem;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:723:7  */
  assign n7658_o = new_i ? n7958_o : n7652_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:723:7  */
  assign n7659_o = new_i ? n8093_o : n7657_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:756:60  */
  assign n7694_o = acc_tag_ff == tag_mem_rd;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:756:44  */
  assign n7695_o = n7694_o & valid_mem_rd;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:756:18  */
  assign n7696_o = n7695_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:757:44  */
  assign n7699_o = dirty_mem_rd & valid_mem_rd;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:757:69  */
  assign n7701_o = 1'b1 & n7699_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:757:18  */
  assign n7702_o = n7701_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:771:15  */
  assign n7707_o = we_i[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:772:62  */
  assign n7712_o = wdata_i[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:774:15  */
  assign n7715_o = we_i[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:775:62  */
  assign n7720_o = wdata_i[15:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:777:15  */
  assign n7723_o = we_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:778:62  */
  assign n7728_o = wdata_i[23:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:780:15  */
  assign n7731_o = we_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:781:62  */
  assign n7736_o = wdata_i[31:24]; // extract
  assign n7770_o = {n7819_data, n7816_data, n7813_data, n7810_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:797:26  */
  assign n7775_o = stat_mem_rd & valid_mem_rd;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:722:5  */
  always @(posedge clk_i or posedge n7638_o)
    if (n7638_o)
      n7776_q <= 32'b00000000000000000000000000000000;
    else
      n7776_q <= n7658_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:722:5  */
  always @(posedge clk_i or posedge n7638_o)
    if (n7638_o)
      n7777_q <= 32'b00000000000000000000000000000000;
    else
      n7777_q <= n7659_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:717:3  */
  assign n7778_o = ~n7638_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:722:5  */
  assign n7779_o = n7778_o ? n8417_o : valid_mem_rd;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:722:5  */
  always @(posedge clk_i)
    n7780_q <= n7779_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:717:3  */
  assign n7781_o = ~n7638_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:722:5  */
  assign n7782_o = n7781_o ? n8471_o : dirty_mem_rd;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:722:5  */
  always @(posedge clk_i)
    n7783_q <= n7782_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:708:5  */
  always @(posedge clk_i or posedge n7628_o)
    if (n7628_o)
      n7799_q <= 22'b0000000000000000000000;
    else
      n7799_q <= acc_tag;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:708:5  */
  always @(posedge clk_i or posedge n7628_o)
    if (n7628_o)
      n7800_q <= 5'b00000;
    else
      n7800_q <= acc_idx;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:705:5  */
  assign n7801_o = {tag_mem_rd, acc_idx_ff, 5'b00000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:749:29  */
  reg [21:0] tag_mem[31:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n7803_data <= tag_mem[acc_idx];
  always @(posedge clk_i)
    if (new_i)
      tag_mem[acc_idx] <= acc_tag;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:749:29  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:747:17  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:787:48  */
  reg [7:0] data_mem_b0[255:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n7810_data <= data_mem_b0[acc_adr];
  always @(posedge clk_i)
    if (n7707_o)
      data_mem_b0[acc_adr] <= n7712_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:675:10  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:772:21  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:788:48  */
  reg [7:0] data_mem_b1[255:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n7813_data <= data_mem_b1[acc_adr];
  always @(posedge clk_i)
    if (n7715_o)
      data_mem_b1[acc_adr] <= n7720_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:788:48  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:775:21  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:789:48  */
  reg [7:0] data_mem_b2[255:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n7816_data <= data_mem_b2[acc_adr];
  always @(posedge clk_i)
    if (n7723_o)
      data_mem_b2[acc_adr] <= n7728_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:789:48  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:778:21  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:790:48  */
  reg [7:0] data_mem_b3[255:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n7819_data <= data_mem_b3[acc_adr];
  always @(posedge clk_i)
    if (n7731_o)
      data_mem_b3[acc_adr] <= n7736_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:790:48  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:781:21  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:680:49  */
  reg stat_mem[255:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n7822_data <= stat_mem[acc_adr];
  always @(posedge clk_i)
    if (swe_i)
      stat_mem[acc_adr] <= wstat_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:769:5  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:784:18  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7824_o = acc_idx[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7825_o = ~n7824_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7826_o = acc_idx[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7827_o = ~n7826_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7828_o = n7825_o & n7827_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7829_o = n7825_o & n7826_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7830_o = n7824_o & n7827_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7831_o = n7824_o & n7826_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7832_o = acc_idx[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7833_o = ~n7832_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7834_o = n7828_o & n7833_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7835_o = n7828_o & n7832_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7836_o = n7829_o & n7833_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7837_o = n7829_o & n7832_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7838_o = n7830_o & n7833_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7839_o = n7830_o & n7832_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7840_o = n7831_o & n7833_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7841_o = n7831_o & n7832_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7842_o = acc_idx[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7843_o = ~n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7844_o = n7834_o & n7843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7845_o = n7834_o & n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7846_o = n7835_o & n7843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7847_o = n7835_o & n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7848_o = n7836_o & n7843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7849_o = n7836_o & n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7850_o = n7837_o & n7843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7851_o = n7837_o & n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7852_o = n7838_o & n7843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7853_o = n7838_o & n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7854_o = n7839_o & n7843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7855_o = n7839_o & n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7856_o = n7840_o & n7843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7857_o = n7840_o & n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7858_o = n7841_o & n7843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7859_o = n7841_o & n7842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7860_o = acc_idx[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7861_o = ~n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7862_o = n7844_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7863_o = n7844_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7864_o = n7845_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7865_o = n7845_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7866_o = n7846_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7867_o = n7846_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7868_o = n7847_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7869_o = n7847_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7870_o = n7848_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7871_o = n7848_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7872_o = n7849_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7873_o = n7849_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7874_o = n7850_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7875_o = n7850_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7876_o = n7851_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7877_o = n7851_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7878_o = n7852_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7879_o = n7852_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7880_o = n7853_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7881_o = n7853_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7882_o = n7854_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7883_o = n7854_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7884_o = n7855_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7885_o = n7855_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7886_o = n7856_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7887_o = n7856_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7888_o = n7857_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7889_o = n7857_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7890_o = n7858_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7891_o = n7858_o & n7860_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7892_o = n7859_o & n7861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7893_o = n7859_o & n7860_o;
  assign n7894_o = valid_mem[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7895_o = n7862_o ? 1'b1 : n7894_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:705:5  */
  assign n7896_o = valid_mem[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7897_o = n7863_o ? 1'b1 : n7896_o;
  assign n7898_o = valid_mem[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7899_o = n7864_o ? 1'b1 : n7898_o;
  assign n7900_o = valid_mem[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7901_o = n7865_o ? 1'b1 : n7900_o;
  assign n7902_o = valid_mem[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7903_o = n7866_o ? 1'b1 : n7902_o;
  assign n7904_o = valid_mem[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7905_o = n7867_o ? 1'b1 : n7904_o;
  assign n7906_o = valid_mem[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7907_o = n7868_o ? 1'b1 : n7906_o;
  assign n7908_o = valid_mem[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7909_o = n7869_o ? 1'b1 : n7908_o;
  assign n7910_o = valid_mem[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7911_o = n7870_o ? 1'b1 : n7910_o;
  assign n7912_o = valid_mem[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7913_o = n7871_o ? 1'b1 : n7912_o;
  assign n7914_o = valid_mem[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7915_o = n7872_o ? 1'b1 : n7914_o;
  assign n7916_o = valid_mem[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7917_o = n7873_o ? 1'b1 : n7916_o;
  assign n7918_o = valid_mem[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7919_o = n7874_o ? 1'b1 : n7918_o;
  assign n7920_o = valid_mem[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7921_o = n7875_o ? 1'b1 : n7920_o;
  assign n7922_o = valid_mem[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7923_o = n7876_o ? 1'b1 : n7922_o;
  assign n7924_o = valid_mem[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7925_o = n7877_o ? 1'b1 : n7924_o;
  assign n7926_o = valid_mem[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7927_o = n7878_o ? 1'b1 : n7926_o;
  assign n7928_o = valid_mem[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7929_o = n7879_o ? 1'b1 : n7928_o;
  assign n7930_o = valid_mem[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7931_o = n7880_o ? 1'b1 : n7930_o;
  assign n7932_o = valid_mem[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7933_o = n7881_o ? 1'b1 : n7932_o;
  assign n7934_o = valid_mem[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7935_o = n7882_o ? 1'b1 : n7934_o;
  assign n7936_o = valid_mem[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7937_o = n7883_o ? 1'b1 : n7936_o;
  assign n7938_o = valid_mem[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7939_o = n7884_o ? 1'b1 : n7938_o;
  assign n7940_o = valid_mem[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7941_o = n7885_o ? 1'b1 : n7940_o;
  assign n7942_o = valid_mem[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7943_o = n7886_o ? 1'b1 : n7942_o;
  assign n7944_o = valid_mem[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7945_o = n7887_o ? 1'b1 : n7944_o;
  assign n7946_o = valid_mem[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7947_o = n7888_o ? 1'b1 : n7946_o;
  assign n7948_o = valid_mem[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7949_o = n7889_o ? 1'b1 : n7948_o;
  assign n7950_o = valid_mem[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7951_o = n7890_o ? 1'b1 : n7950_o;
  assign n7952_o = valid_mem[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7953_o = n7891_o ? 1'b1 : n7952_o;
  assign n7954_o = valid_mem[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7955_o = n7892_o ? 1'b1 : n7954_o;
  assign n7956_o = valid_mem[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:724:9  */
  assign n7957_o = n7893_o ? 1'b1 : n7956_o;
  assign n7958_o = {n7957_o, n7955_o, n7953_o, n7951_o, n7949_o, n7947_o, n7945_o, n7943_o, n7941_o, n7939_o, n7937_o, n7935_o, n7933_o, n7931_o, n7929_o, n7927_o, n7925_o, n7923_o, n7921_o, n7919_o, n7917_o, n7915_o, n7913_o, n7911_o, n7909_o, n7907_o, n7905_o, n7903_o, n7901_o, n7899_o, n7897_o, n7895_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7959_o = acc_idx[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7960_o = ~n7959_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7961_o = acc_idx[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7962_o = ~n7961_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7963_o = n7960_o & n7962_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7964_o = n7960_o & n7961_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7965_o = n7959_o & n7962_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7966_o = n7959_o & n7961_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7967_o = acc_idx[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7968_o = ~n7967_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7969_o = n7963_o & n7968_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7970_o = n7963_o & n7967_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7971_o = n7964_o & n7968_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7972_o = n7964_o & n7967_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7973_o = n7965_o & n7968_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7974_o = n7965_o & n7967_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7975_o = n7966_o & n7968_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7976_o = n7966_o & n7967_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7977_o = acc_idx[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7978_o = ~n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7979_o = n7969_o & n7978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7980_o = n7969_o & n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7981_o = n7970_o & n7978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7982_o = n7970_o & n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7983_o = n7971_o & n7978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7984_o = n7971_o & n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7985_o = n7972_o & n7978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7986_o = n7972_o & n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7987_o = n7973_o & n7978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7988_o = n7973_o & n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7989_o = n7974_o & n7978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7990_o = n7974_o & n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7991_o = n7975_o & n7978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7992_o = n7975_o & n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7993_o = n7976_o & n7978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7994_o = n7976_o & n7977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7995_o = acc_idx[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7996_o = ~n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7997_o = n7979_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7998_o = n7979_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n7999_o = n7980_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8000_o = n7980_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8001_o = n7981_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8002_o = n7981_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8003_o = n7982_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8004_o = n7982_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8005_o = n7983_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8006_o = n7983_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8007_o = n7984_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8008_o = n7984_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8009_o = n7985_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8010_o = n7985_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8011_o = n7986_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8012_o = n7986_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8013_o = n7987_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8014_o = n7987_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8015_o = n7988_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8016_o = n7988_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8017_o = n7989_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8018_o = n7989_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8019_o = n7990_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8020_o = n7990_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8021_o = n7991_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8022_o = n7991_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8023_o = n7992_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8024_o = n7992_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8025_o = n7993_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8026_o = n7993_o & n7995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8027_o = n7994_o & n7996_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8028_o = n7994_o & n7995_o;
  assign n8029_o = dirty_mem[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8030_o = n7997_o ? 1'b0 : n8029_o;
  assign n8031_o = dirty_mem[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8032_o = n7998_o ? 1'b0 : n8031_o;
  assign n8033_o = dirty_mem[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8034_o = n7999_o ? 1'b0 : n8033_o;
  assign n8035_o = dirty_mem[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8036_o = n8000_o ? 1'b0 : n8035_o;
  assign n8037_o = dirty_mem[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8038_o = n8001_o ? 1'b0 : n8037_o;
  assign n8039_o = dirty_mem[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8040_o = n8002_o ? 1'b0 : n8039_o;
  assign n8041_o = dirty_mem[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8042_o = n8003_o ? 1'b0 : n8041_o;
  assign n8043_o = dirty_mem[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8044_o = n8004_o ? 1'b0 : n8043_o;
  assign n8045_o = dirty_mem[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8046_o = n8005_o ? 1'b0 : n8045_o;
  assign n8047_o = dirty_mem[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8048_o = n8006_o ? 1'b0 : n8047_o;
  assign n8049_o = dirty_mem[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8050_o = n8007_o ? 1'b0 : n8049_o;
  assign n8051_o = dirty_mem[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8052_o = n8008_o ? 1'b0 : n8051_o;
  assign n8053_o = dirty_mem[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8054_o = n8009_o ? 1'b0 : n8053_o;
  assign n8055_o = dirty_mem[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8056_o = n8010_o ? 1'b0 : n8055_o;
  assign n8057_o = dirty_mem[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8058_o = n8011_o ? 1'b0 : n8057_o;
  assign n8059_o = dirty_mem[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8060_o = n8012_o ? 1'b0 : n8059_o;
  assign n8061_o = dirty_mem[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8062_o = n8013_o ? 1'b0 : n8061_o;
  assign n8063_o = dirty_mem[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8064_o = n8014_o ? 1'b0 : n8063_o;
  assign n8065_o = dirty_mem[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8066_o = n8015_o ? 1'b0 : n8065_o;
  assign n8067_o = dirty_mem[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8068_o = n8016_o ? 1'b0 : n8067_o;
  assign n8069_o = dirty_mem[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8070_o = n8017_o ? 1'b0 : n8069_o;
  assign n8071_o = dirty_mem[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8072_o = n8018_o ? 1'b0 : n8071_o;
  assign n8073_o = dirty_mem[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8074_o = n8019_o ? 1'b0 : n8073_o;
  assign n8075_o = dirty_mem[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8076_o = n8020_o ? 1'b0 : n8075_o;
  assign n8077_o = dirty_mem[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8078_o = n8021_o ? 1'b0 : n8077_o;
  assign n8079_o = dirty_mem[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8080_o = n8022_o ? 1'b0 : n8079_o;
  assign n8081_o = dirty_mem[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8082_o = n8023_o ? 1'b0 : n8081_o;
  assign n8083_o = dirty_mem[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8084_o = n8024_o ? 1'b0 : n8083_o;
  assign n8085_o = dirty_mem[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8086_o = n8025_o ? 1'b0 : n8085_o;
  assign n8087_o = dirty_mem[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8088_o = n8026_o ? 1'b0 : n8087_o;
  assign n8089_o = dirty_mem[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8090_o = n8027_o ? 1'b0 : n8089_o;
  assign n8091_o = dirty_mem[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:725:9  */
  assign n8092_o = n8028_o ? 1'b0 : n8091_o;
  assign n8093_o = {n8092_o, n8090_o, n8088_o, n8086_o, n8084_o, n8082_o, n8080_o, n8078_o, n8076_o, n8074_o, n8072_o, n8070_o, n8068_o, n8066_o, n8064_o, n8062_o, n8060_o, n8058_o, n8056_o, n8054_o, n8052_o, n8050_o, n8048_o, n8046_o, n8044_o, n8042_o, n8040_o, n8038_o, n8036_o, n8034_o, n8032_o, n8030_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8094_o = acc_idx[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8095_o = ~n8094_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8096_o = acc_idx[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8097_o = ~n8096_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8098_o = n8095_o & n8097_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8099_o = n8095_o & n8096_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8100_o = n8094_o & n8097_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8101_o = n8094_o & n8096_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8102_o = acc_idx[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8103_o = ~n8102_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8104_o = n8098_o & n8103_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8105_o = n8098_o & n8102_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8106_o = n8099_o & n8103_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8107_o = n8099_o & n8102_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8108_o = n8100_o & n8103_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8109_o = n8100_o & n8102_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8110_o = n8101_o & n8103_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8111_o = n8101_o & n8102_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8112_o = acc_idx[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8113_o = ~n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8114_o = n8104_o & n8113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8115_o = n8104_o & n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8116_o = n8105_o & n8113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8117_o = n8105_o & n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8118_o = n8106_o & n8113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8119_o = n8106_o & n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8120_o = n8107_o & n8113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8121_o = n8107_o & n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8122_o = n8108_o & n8113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8123_o = n8108_o & n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8124_o = n8109_o & n8113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8125_o = n8109_o & n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8126_o = n8110_o & n8113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8127_o = n8110_o & n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8128_o = n8111_o & n8113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8129_o = n8111_o & n8112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8130_o = acc_idx[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8131_o = ~n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8132_o = n8114_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8133_o = n8114_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8134_o = n8115_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8135_o = n8115_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8136_o = n8116_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8137_o = n8116_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8138_o = n8117_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8139_o = n8117_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8140_o = n8118_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8141_o = n8118_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8142_o = n8119_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8143_o = n8119_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8144_o = n8120_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8145_o = n8120_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8146_o = n8121_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8147_o = n8121_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8148_o = n8122_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8149_o = n8122_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8150_o = n8123_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8151_o = n8123_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8152_o = n8124_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8153_o = n8124_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8154_o = n8125_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8155_o = n8125_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8156_o = n8126_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8157_o = n8126_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8158_o = n8127_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8159_o = n8127_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8160_o = n8128_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8161_o = n8128_o & n8130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8162_o = n8129_o & n8131_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8163_o = n8129_o & n8130_o;
  assign n8164_o = valid_mem[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8165_o = n8132_o ? 1'b0 : n8164_o;
  assign n8166_o = valid_mem[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8167_o = n8133_o ? 1'b0 : n8166_o;
  assign n8168_o = valid_mem[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8169_o = n8134_o ? 1'b0 : n8168_o;
  assign n8170_o = valid_mem[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8171_o = n8135_o ? 1'b0 : n8170_o;
  assign n8172_o = valid_mem[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8173_o = n8136_o ? 1'b0 : n8172_o;
  assign n8174_o = valid_mem[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8175_o = n8137_o ? 1'b0 : n8174_o;
  assign n8176_o = valid_mem[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8177_o = n8138_o ? 1'b0 : n8176_o;
  assign n8178_o = valid_mem[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8179_o = n8139_o ? 1'b0 : n8178_o;
  assign n8180_o = valid_mem[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8181_o = n8140_o ? 1'b0 : n8180_o;
  assign n8182_o = valid_mem[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8183_o = n8141_o ? 1'b0 : n8182_o;
  assign n8184_o = valid_mem[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8185_o = n8142_o ? 1'b0 : n8184_o;
  assign n8186_o = valid_mem[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8187_o = n8143_o ? 1'b0 : n8186_o;
  assign n8188_o = valid_mem[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8189_o = n8144_o ? 1'b0 : n8188_o;
  assign n8190_o = valid_mem[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8191_o = n8145_o ? 1'b0 : n8190_o;
  assign n8192_o = valid_mem[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8193_o = n8146_o ? 1'b0 : n8192_o;
  assign n8194_o = valid_mem[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8195_o = n8147_o ? 1'b0 : n8194_o;
  assign n8196_o = valid_mem[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8197_o = n8148_o ? 1'b0 : n8196_o;
  assign n8198_o = valid_mem[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8199_o = n8149_o ? 1'b0 : n8198_o;
  assign n8200_o = valid_mem[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8201_o = n8150_o ? 1'b0 : n8200_o;
  assign n8202_o = valid_mem[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8203_o = n8151_o ? 1'b0 : n8202_o;
  assign n8204_o = valid_mem[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8205_o = n8152_o ? 1'b0 : n8204_o;
  assign n8206_o = valid_mem[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8207_o = n8153_o ? 1'b0 : n8206_o;
  assign n8208_o = valid_mem[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8209_o = n8154_o ? 1'b0 : n8208_o;
  assign n8210_o = valid_mem[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8211_o = n8155_o ? 1'b0 : n8210_o;
  assign n8212_o = valid_mem[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8213_o = n8156_o ? 1'b0 : n8212_o;
  assign n8214_o = valid_mem[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8215_o = n8157_o ? 1'b0 : n8214_o;
  assign n8216_o = valid_mem[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8217_o = n8158_o ? 1'b0 : n8216_o;
  assign n8218_o = valid_mem[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8219_o = n8159_o ? 1'b0 : n8218_o;
  assign n8220_o = valid_mem[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8221_o = n8160_o ? 1'b0 : n8220_o;
  assign n8222_o = valid_mem[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8223_o = n8161_o ? 1'b0 : n8222_o;
  assign n8224_o = valid_mem[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8225_o = n8162_o ? 1'b0 : n8224_o;
  assign n8226_o = valid_mem[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:728:11  */
  assign n8227_o = n8163_o ? 1'b0 : n8226_o;
  assign n8228_o = {n8227_o, n8225_o, n8223_o, n8221_o, n8219_o, n8217_o, n8215_o, n8213_o, n8211_o, n8209_o, n8207_o, n8205_o, n8203_o, n8201_o, n8199_o, n8197_o, n8195_o, n8193_o, n8191_o, n8189_o, n8187_o, n8185_o, n8183_o, n8181_o, n8179_o, n8177_o, n8175_o, n8173_o, n8171_o, n8169_o, n8167_o, n8165_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8229_o = acc_idx[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8230_o = ~n8229_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8231_o = acc_idx[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8232_o = ~n8231_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8233_o = n8230_o & n8232_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8234_o = n8230_o & n8231_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8235_o = n8229_o & n8232_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8236_o = n8229_o & n8231_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8237_o = acc_idx[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8238_o = ~n8237_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8239_o = n8233_o & n8238_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8240_o = n8233_o & n8237_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8241_o = n8234_o & n8238_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8242_o = n8234_o & n8237_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8243_o = n8235_o & n8238_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8244_o = n8235_o & n8237_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8245_o = n8236_o & n8238_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8246_o = n8236_o & n8237_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8247_o = acc_idx[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8248_o = ~n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8249_o = n8239_o & n8248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8250_o = n8239_o & n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8251_o = n8240_o & n8248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8252_o = n8240_o & n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8253_o = n8241_o & n8248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8254_o = n8241_o & n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8255_o = n8242_o & n8248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8256_o = n8242_o & n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8257_o = n8243_o & n8248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8258_o = n8243_o & n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8259_o = n8244_o & n8248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8260_o = n8244_o & n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8261_o = n8245_o & n8248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8262_o = n8245_o & n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8263_o = n8246_o & n8248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8264_o = n8246_o & n8247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8265_o = acc_idx[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8266_o = ~n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8267_o = n8249_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8268_o = n8249_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8269_o = n8250_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8270_o = n8250_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8271_o = n8251_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8272_o = n8251_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8273_o = n8252_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8274_o = n8252_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8275_o = n8253_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8276_o = n8253_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8277_o = n8254_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8278_o = n8254_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8279_o = n8255_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8280_o = n8255_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8281_o = n8256_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8282_o = n8256_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8283_o = n8257_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8284_o = n8257_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8285_o = n8258_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8286_o = n8258_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8287_o = n8259_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8288_o = n8259_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8289_o = n8260_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8290_o = n8260_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8291_o = n8261_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8292_o = n8261_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8293_o = n8262_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8294_o = n8262_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8295_o = n8263_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8296_o = n8263_o & n8265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8297_o = n8264_o & n8266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8298_o = n8264_o & n8265_o;
  assign n8299_o = dirty_mem[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8300_o = n8267_o ? 1'b1 : n8299_o;
  assign n8301_o = dirty_mem[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8302_o = n8268_o ? 1'b1 : n8301_o;
  assign n8303_o = dirty_mem[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8304_o = n8269_o ? 1'b1 : n8303_o;
  assign n8305_o = dirty_mem[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8306_o = n8270_o ? 1'b1 : n8305_o;
  assign n8307_o = dirty_mem[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8308_o = n8271_o ? 1'b1 : n8307_o;
  assign n8309_o = dirty_mem[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8310_o = n8272_o ? 1'b1 : n8309_o;
  assign n8311_o = dirty_mem[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8312_o = n8273_o ? 1'b1 : n8311_o;
  assign n8313_o = dirty_mem[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8314_o = n8274_o ? 1'b1 : n8313_o;
  assign n8315_o = dirty_mem[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8316_o = n8275_o ? 1'b1 : n8315_o;
  assign n8317_o = dirty_mem[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8318_o = n8276_o ? 1'b1 : n8317_o;
  assign n8319_o = dirty_mem[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8320_o = n8277_o ? 1'b1 : n8319_o;
  assign n8321_o = dirty_mem[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8322_o = n8278_o ? 1'b1 : n8321_o;
  assign n8323_o = dirty_mem[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8324_o = n8279_o ? 1'b1 : n8323_o;
  assign n8325_o = dirty_mem[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8326_o = n8280_o ? 1'b1 : n8325_o;
  assign n8327_o = dirty_mem[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8328_o = n8281_o ? 1'b1 : n8327_o;
  assign n8329_o = dirty_mem[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8330_o = n8282_o ? 1'b1 : n8329_o;
  assign n8331_o = dirty_mem[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8332_o = n8283_o ? 1'b1 : n8331_o;
  assign n8333_o = dirty_mem[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8334_o = n8284_o ? 1'b1 : n8333_o;
  assign n8335_o = dirty_mem[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8336_o = n8285_o ? 1'b1 : n8335_o;
  assign n8337_o = dirty_mem[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8338_o = n8286_o ? 1'b1 : n8337_o;
  assign n8339_o = dirty_mem[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8340_o = n8287_o ? 1'b1 : n8339_o;
  assign n8341_o = dirty_mem[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8342_o = n8288_o ? 1'b1 : n8341_o;
  assign n8343_o = dirty_mem[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8344_o = n8289_o ? 1'b1 : n8343_o;
  assign n8345_o = dirty_mem[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8346_o = n8290_o ? 1'b1 : n8345_o;
  assign n8347_o = dirty_mem[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8348_o = n8291_o ? 1'b1 : n8347_o;
  assign n8349_o = dirty_mem[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8350_o = n8292_o ? 1'b1 : n8349_o;
  assign n8351_o = dirty_mem[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8352_o = n8293_o ? 1'b1 : n8351_o;
  assign n8353_o = dirty_mem[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8354_o = n8294_o ? 1'b1 : n8353_o;
  assign n8355_o = dirty_mem[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8356_o = n8295_o ? 1'b1 : n8355_o;
  assign n8357_o = dirty_mem[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8358_o = n8296_o ? 1'b1 : n8357_o;
  assign n8359_o = dirty_mem[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8360_o = n8297_o ? 1'b1 : n8359_o;
  assign n8361_o = dirty_mem[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8362_o = n8298_o ? 1'b1 : n8361_o;
  assign n8363_o = {n8362_o, n8360_o, n8358_o, n8356_o, n8354_o, n8352_o, n8350_o, n8348_o, n8346_o, n8344_o, n8342_o, n8340_o, n8338_o, n8336_o, n8334_o, n8332_o, n8330_o, n8328_o, n8326_o, n8324_o, n8322_o, n8320_o, n8318_o, n8316_o, n8314_o, n8312_o, n8310_o, n8308_o, n8306_o, n8304_o, n8302_o, n8300_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:21  */
  assign n8364_o = valid_mem[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:731:11  */
  assign n8365_o = valid_mem[1]; // extract
  assign n8366_o = valid_mem[2]; // extract
  assign n8367_o = valid_mem[3]; // extract
  assign n8368_o = valid_mem[4]; // extract
  assign n8369_o = valid_mem[5]; // extract
  assign n8370_o = valid_mem[6]; // extract
  assign n8371_o = valid_mem[7]; // extract
  assign n8372_o = valid_mem[8]; // extract
  assign n8373_o = valid_mem[9]; // extract
  assign n8374_o = valid_mem[10]; // extract
  assign n8375_o = valid_mem[11]; // extract
  assign n8376_o = valid_mem[12]; // extract
  assign n8377_o = valid_mem[13]; // extract
  assign n8378_o = valid_mem[14]; // extract
  assign n8379_o = valid_mem[15]; // extract
  assign n8380_o = valid_mem[16]; // extract
  assign n8381_o = valid_mem[17]; // extract
  assign n8382_o = valid_mem[18]; // extract
  assign n8383_o = valid_mem[19]; // extract
  assign n8384_o = valid_mem[20]; // extract
  assign n8385_o = valid_mem[21]; // extract
  assign n8386_o = valid_mem[22]; // extract
  assign n8387_o = valid_mem[23]; // extract
  assign n8388_o = valid_mem[24]; // extract
  assign n8389_o = valid_mem[25]; // extract
  assign n8390_o = valid_mem[26]; // extract
  assign n8391_o = valid_mem[27]; // extract
  assign n8392_o = valid_mem[28]; // extract
  assign n8393_o = valid_mem[29]; // extract
  assign n8394_o = valid_mem[30]; // extract
  assign n8395_o = valid_mem[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8396_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8396_o)
      2'b00: n8397_o = n8364_o;
      2'b01: n8397_o = n8365_o;
      2'b10: n8397_o = n8366_o;
      2'b11: n8397_o = n8367_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8398_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8398_o)
      2'b00: n8399_o = n8368_o;
      2'b01: n8399_o = n8369_o;
      2'b10: n8399_o = n8370_o;
      2'b11: n8399_o = n8371_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8400_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8400_o)
      2'b00: n8401_o = n8372_o;
      2'b01: n8401_o = n8373_o;
      2'b10: n8401_o = n8374_o;
      2'b11: n8401_o = n8375_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8402_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8402_o)
      2'b00: n8403_o = n8376_o;
      2'b01: n8403_o = n8377_o;
      2'b10: n8403_o = n8378_o;
      2'b11: n8403_o = n8379_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8404_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8404_o)
      2'b00: n8405_o = n8380_o;
      2'b01: n8405_o = n8381_o;
      2'b10: n8405_o = n8382_o;
      2'b11: n8405_o = n8383_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8406_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8406_o)
      2'b00: n8407_o = n8384_o;
      2'b01: n8407_o = n8385_o;
      2'b10: n8407_o = n8386_o;
      2'b11: n8407_o = n8387_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8408_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8408_o)
      2'b00: n8409_o = n8388_o;
      2'b01: n8409_o = n8389_o;
      2'b10: n8409_o = n8390_o;
      2'b11: n8409_o = n8391_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8410_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8410_o)
      2'b00: n8411_o = n8392_o;
      2'b01: n8411_o = n8393_o;
      2'b10: n8411_o = n8394_o;
      2'b11: n8411_o = n8395_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8412_o = acc_idx[3:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8412_o)
      2'b00: n8413_o = n8397_o;
      2'b01: n8413_o = n8399_o;
      2'b10: n8413_o = n8401_o;
      2'b11: n8413_o = n8403_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8414_o = acc_idx[3:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  always @*
    case (n8414_o)
      2'b00: n8415_o = n8405_o;
      2'b01: n8415_o = n8407_o;
      2'b10: n8415_o = n8409_o;
      2'b11: n8415_o = n8411_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8416_o = acc_idx[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8417_o = n8416_o ? n8415_o : n8413_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:32  */
  assign n8418_o = dirty_mem[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:735:33  */
  assign n8419_o = dirty_mem[1]; // extract
  assign n8420_o = dirty_mem[2]; // extract
  assign n8421_o = dirty_mem[3]; // extract
  assign n8422_o = dirty_mem[4]; // extract
  assign n8423_o = dirty_mem[5]; // extract
  assign n8424_o = dirty_mem[6]; // extract
  assign n8425_o = dirty_mem[7]; // extract
  assign n8426_o = dirty_mem[8]; // extract
  assign n8427_o = dirty_mem[9]; // extract
  assign n8428_o = dirty_mem[10]; // extract
  assign n8429_o = dirty_mem[11]; // extract
  assign n8430_o = dirty_mem[12]; // extract
  assign n8431_o = dirty_mem[13]; // extract
  assign n8432_o = dirty_mem[14]; // extract
  assign n8433_o = dirty_mem[15]; // extract
  assign n8434_o = dirty_mem[16]; // extract
  assign n8435_o = dirty_mem[17]; // extract
  assign n8436_o = dirty_mem[18]; // extract
  assign n8437_o = dirty_mem[19]; // extract
  assign n8438_o = dirty_mem[20]; // extract
  assign n8439_o = dirty_mem[21]; // extract
  assign n8440_o = dirty_mem[22]; // extract
  assign n8441_o = dirty_mem[23]; // extract
  assign n8442_o = dirty_mem[24]; // extract
  assign n8443_o = dirty_mem[25]; // extract
  assign n8444_o = dirty_mem[26]; // extract
  assign n8445_o = dirty_mem[27]; // extract
  assign n8446_o = dirty_mem[28]; // extract
  assign n8447_o = dirty_mem[29]; // extract
  assign n8448_o = dirty_mem[30]; // extract
  assign n8449_o = dirty_mem[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8450_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8450_o)
      2'b00: n8451_o = n8418_o;
      2'b01: n8451_o = n8419_o;
      2'b10: n8451_o = n8420_o;
      2'b11: n8451_o = n8421_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8452_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8452_o)
      2'b00: n8453_o = n8422_o;
      2'b01: n8453_o = n8423_o;
      2'b10: n8453_o = n8424_o;
      2'b11: n8453_o = n8425_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8454_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8454_o)
      2'b00: n8455_o = n8426_o;
      2'b01: n8455_o = n8427_o;
      2'b10: n8455_o = n8428_o;
      2'b11: n8455_o = n8429_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8456_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8456_o)
      2'b00: n8457_o = n8430_o;
      2'b01: n8457_o = n8431_o;
      2'b10: n8457_o = n8432_o;
      2'b11: n8457_o = n8433_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8458_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8458_o)
      2'b00: n8459_o = n8434_o;
      2'b01: n8459_o = n8435_o;
      2'b10: n8459_o = n8436_o;
      2'b11: n8459_o = n8437_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8460_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8460_o)
      2'b00: n8461_o = n8438_o;
      2'b01: n8461_o = n8439_o;
      2'b10: n8461_o = n8440_o;
      2'b11: n8461_o = n8441_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8462_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8462_o)
      2'b00: n8463_o = n8442_o;
      2'b01: n8463_o = n8443_o;
      2'b10: n8463_o = n8444_o;
      2'b11: n8463_o = n8445_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8464_o = acc_idx[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8464_o)
      2'b00: n8465_o = n8446_o;
      2'b01: n8465_o = n8447_o;
      2'b10: n8465_o = n8448_o;
      2'b11: n8465_o = n8449_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8466_o = acc_idx[3:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8466_o)
      2'b00: n8467_o = n8451_o;
      2'b01: n8467_o = n8453_o;
      2'b10: n8467_o = n8455_o;
      2'b11: n8467_o = n8457_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8468_o = acc_idx[3:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  always @*
    case (n8468_o)
      2'b00: n8469_o = n8459_o;
      2'b01: n8469_o = n8461_o;
      2'b10: n8469_o = n8463_o;
      2'b11: n8469_o = n8465_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8470_o = acc_idx[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:736:32  */
  assign n8471_o = n8470_o ? n8469_o : n8467_o;
endmodule

module neorv32_cache_host_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  rstn_i,
   input  clk_i,
   input  [31:0] req_i_addr,
   input  [31:0] req_i_data,
   input  [3:0] req_i_ben,
   input  req_i_stb,
   input  req_i_rw,
   input  req_i_src,
   input  req_i_priv,
   input  req_i_rvso,
   input  req_i_fence,
   input  bus_busy_i,
   input  hit_i,
   input  [31:0] rdata_i,
   input  rstat_i,
   output [31:0] rsp_o_data,
   output rsp_o_ack,
   output rsp_o_err,
   output bus_sync_o,
   output bus_miss_o,
   output dirty_o,
   output [31:0] addr_o,
   output [3:0] we_o,
   output swe_o,
   output [31:0] wdata_o,
   output wstat_o);
  wire [73:0] n7484_o;
  wire [31:0] n7486_o;
  wire n7487_o;
  wire n7488_o;
  wire [9:0] ctrl;
  wire n7498_o;
  wire [2:0] n7503_o;
  wire n7504_o;
  wire n7505_o;
  wire [2:0] n7517_o;
  wire n7518_o;
  wire n7519_o;
  wire n7520_o;
  wire n7521_o;
  wire n7522_o;
  wire n7523_o;
  wire [31:0] n7524_o;
  wire [31:0] n7525_o;
  wire [2:0] n7526_o;
  wire n7527_o;
  wire n7529_o;
  wire n7530_o;
  wire n7531_o;
  wire [2:0] n7534_o;
  wire n7537_o;
  wire [2:0] n7538_o;
  wire n7540_o;
  wire n7542_o;
  wire n7544_o;
  wire [3:0] n7545_o;
  wire n7548_o;
  wire [3:0] n7550_o;
  wire n7551_o;
  wire [1:0] n7554_o;
  wire [1:0] n7556_o;
  wire n7559_o;
  wire n7561_o;
  wire [3:0] n7563_o;
  wire [2:0] n7564_o;
  wire n7566_o;
  wire n7568_o;
  wire [2:0] n7570_o;
  wire n7572_o;
  wire n7573_o;
  wire [2:0] n7575_o;
  wire n7577_o;
  wire n7581_o;
  wire [4:0] n7583_o;
  reg [31:0] n7585_o;
  wire n7586_o;
  reg n7588_o;
  wire n7589_o;
  reg n7591_o;
  reg n7596_o;
  reg n7599_o;
  reg n7602_o;
  reg [3:0] n7605_o;
  reg [2:0] n7607_o;
  reg n7608_o;
  reg n7609_o;
  localparam n7611_o = 1'b0;
  localparam n7612_o = 1'b0;
  reg n7613_q;
  reg n7614_q;
  reg [2:0] n7615_q;
  wire [9:0] n7616_o;
  wire [33:0] n7617_o;
  assign rsp_o_data = n7486_o; //(module output)
  assign rsp_o_ack = n7487_o; //(module output)
  assign rsp_o_err = n7488_o; //(module output)
  assign bus_sync_o = n7596_o; //(module output)
  assign bus_miss_o = n7599_o; //(module output)
  assign dirty_o = n7602_o; //(module output)
  assign addr_o = n7524_o; //(module output)
  assign we_o = n7605_o; //(module output)
  assign swe_o = n7611_o; //(module output)
  assign wdata_o = n7525_o; //(module output)
  assign wstat_o = n7612_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7484_o = {req_i_fence, req_i_rvso, req_i_priv, req_i_src, req_i_rw, req_i_stb, req_i_ben, req_i_data, req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:133:3  */
  assign n7486_o = n7617_o[31:0]; // extract
  assign n7487_o = n7617_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:108:5  */
  assign n7488_o = n7617_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:483:10  */
  assign ctrl = n7616_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:491:16  */
  assign n7498_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:496:29  */
  assign n7503_o = ctrl[5:3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:497:29  */
  assign n7504_o = ctrl[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:498:29  */
  assign n7505_o = ctrl[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:508:31  */
  assign n7517_o = ctrl[2:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:509:31  */
  assign n7518_o = ctrl[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:509:48  */
  assign n7519_o = n7484_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:509:39  */
  assign n7520_o = n7518_o | n7519_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:510:31  */
  assign n7521_o = ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:510:49  */
  assign n7522_o = n7484_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:510:40  */
  assign n7523_o = n7521_o | n7522_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:514:22  */
  assign n7524_o = n7484_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:517:22  */
  assign n7525_o = n7484_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:15  */
  assign n7526_o = ctrl[2:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:532:18  */
  assign n7527_o = ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:535:22  */
  assign n7529_o = n7484_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:535:42  */
  assign n7530_o = ctrl[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:535:33  */
  assign n7531_o = n7529_o | n7530_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:535:9  */
  assign n7534_o = n7531_o ? 3'b001 : n7517_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:532:9  */
  assign n7537_o = n7527_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:532:9  */
  assign n7538_o = n7527_o ? 3'b011 : n7534_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:530:7  */
  assign n7540_o = n7526_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:548:21  */
  assign n7542_o = n7484_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:548:31  */
  assign n7544_o = 1'b1 & n7542_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:550:30  */
  assign n7545_o = n7484_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:548:11  */
  assign n7548_o = n7544_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:548:11  */
  assign n7550_o = n7544_o ? n7545_o : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:552:29  */
  assign n7551_o = ~rstat_i;
  assign n7554_o = {rstat_i, n7551_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:547:9  */
  assign n7556_o = hit_i ? n7554_o : 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:547:9  */
  assign n7559_o = hit_i ? 1'b0 : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:547:9  */
  assign n7561_o = hit_i ? n7548_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:547:9  */
  assign n7563_o = hit_i ? n7550_o : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:547:9  */
  assign n7564_o = hit_i ? 3'b000 : 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:543:7  */
  assign n7566_o = n7526_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:563:24  */
  assign n7568_o = ~bus_busy_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:563:9  */
  assign n7570_o = n7568_o ? 3'b000 : n7517_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:560:7  */
  assign n7572_o = n7526_o == 3'b011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:569:24  */
  assign n7573_o = ~bus_busy_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:569:9  */
  assign n7575_o = n7573_o ? 3'b001 : n7517_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:567:7  */
  assign n7577_o = n7526_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:573:7  */
  assign n7581_o = n7526_o == 3'b100;
  assign n7583_o = {n7581_o, n7577_o, n7572_o, n7566_o, n7540_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7585_o = 32'b00000000000000000000000000000000;
      5'b01000: n7585_o = 32'b00000000000000000000000000000000;
      5'b00100: n7585_o = 32'b00000000000000000000000000000000;
      5'b00010: n7585_o = rdata_i;
      5'b00001: n7585_o = 32'b00000000000000000000000000000000;
      default: n7585_o = 32'b00000000000000000000000000000000;
    endcase
  assign n7586_o = n7556_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7588_o = 1'b0;
      5'b01000: n7588_o = 1'b0;
      5'b00100: n7588_o = 1'b0;
      5'b00010: n7588_o = n7586_o;
      5'b00001: n7588_o = 1'b0;
      default: n7588_o = 1'b0;
    endcase
  assign n7589_o = n7556_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7591_o = 1'b1;
      5'b01000: n7591_o = 1'b0;
      5'b00100: n7591_o = 1'b0;
      5'b00010: n7591_o = n7589_o;
      5'b00001: n7591_o = 1'b0;
      default: n7591_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7596_o = 1'b0;
      5'b01000: n7596_o = 1'b0;
      5'b00100: n7596_o = 1'b0;
      5'b00010: n7596_o = 1'b0;
      5'b00001: n7596_o = n7537_o;
      default: n7596_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7599_o = 1'b0;
      5'b01000: n7599_o = 1'b0;
      5'b00100: n7599_o = 1'b0;
      5'b00010: n7599_o = n7559_o;
      5'b00001: n7599_o = 1'b0;
      default: n7599_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7602_o = 1'b0;
      5'b01000: n7602_o = 1'b0;
      5'b00100: n7602_o = 1'b0;
      5'b00010: n7602_o = n7561_o;
      5'b00001: n7602_o = 1'b0;
      default: n7602_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7605_o = 4'b0000;
      5'b01000: n7605_o = 4'b0000;
      5'b00100: n7605_o = 4'b0000;
      5'b00010: n7605_o = n7563_o;
      5'b00001: n7605_o = 4'b0000;
      default: n7605_o = 4'b0000;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7607_o = 3'b000;
      5'b01000: n7607_o = n7575_o;
      5'b00100: n7607_o = n7570_o;
      5'b00010: n7607_o = n7564_o;
      5'b00001: n7607_o = n7538_o;
      default: n7607_o = 3'b000;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7608_o = n7520_o;
      5'b01000: n7608_o = n7520_o;
      5'b00100: n7608_o = n7520_o;
      5'b00010: n7608_o = 1'b0;
      5'b00001: n7608_o = n7520_o;
      default: n7608_o = n7520_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:528:5  */
  always @*
    case (n7583_o)
      5'b10000: n7609_o = n7523_o;
      5'b01000: n7609_o = n7523_o;
      5'b00100: n7609_o = 1'b0;
      5'b00010: n7609_o = n7523_o;
      5'b00001: n7609_o = n7523_o;
      default: n7609_o = n7523_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:495:5  */
  always @(posedge clk_i or posedge n7498_o)
    if (n7498_o)
      n7613_q <= 1'b0;
    else
      n7613_q <= n7505_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:495:5  */
  always @(posedge clk_i or posedge n7498_o)
    if (n7498_o)
      n7614_q <= 1'b0;
    else
      n7614_q <= n7504_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:495:5  */
  always @(posedge clk_i or posedge n7498_o)
    if (n7498_o)
      n7615_q <= 3'b000;
    else
      n7615_q <= n7503_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:491:5  */
  assign n7616_o = {n7609_o, n7613_q, n7608_o, n7614_q, n7607_o, n7615_q};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:491:5  */
  assign n7617_o = {n7591_o, n7588_o, n7585_o};
endmodule

module neorv32_cpu_lsu_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_lsu_req,
   input  ctrl_i_lsu_rw,
   input  ctrl_i_lsu_mo_we,
   input  ctrl_i_lsu_fence,
   input  ctrl_i_lsu_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  [31:0] addr_i,
   input  [31:0] wdata_i,
   input  pmp_fault_i,
   input  [31:0] bus_rsp_i_data,
   input  bus_rsp_i_ack,
   input  bus_rsp_i_err,
   output [31:0] rdata_o,
   output [31:0] mar_o,
   output wait_o,
   output ma_load_o,
   output ma_store_o,
   output be_load_o,
   output be_store_o,
   output [31:0] bus_req_o_addr,
   output [31:0] bus_req_o_data,
   output [3:0] bus_req_o_ben,
   output bus_req_o_stb,
   output bus_req_o_rw,
   output bus_req_o_src,
   output bus_req_o_priv,
   output bus_req_o_rvso,
   output bus_req_o_fence);
  wire [66:0] n6687_o;
  wire [31:0] n6696_o;
  wire [31:0] n6697_o;
  wire [3:0] n6698_o;
  wire n6699_o;
  wire n6700_o;
  wire n6701_o;
  wire n6702_o;
  wire n6703_o;
  wire n6704_o;
  wire [33:0] n6705_o;
  wire [31:0] mar;
  wire misaligned;
  wire arbiter_req;
  wire arbiter_err;
  wire n6707_o;
  wire n6709_o;
  wire [1:0] n6710_o;
  wire n6712_o;
  wire n6713_o;
  wire n6715_o;
  wire n6716_o;
  wire n6717_o;
  wire n6718_o;
  wire [1:0] n6719_o;
  reg n6721_o;
  wire n6732_o;
  wire n6737_o;
  wire n6738_o;
  wire n6739_o;
  wire [1:0] n6741_o;
  wire [1:0] n6750_o;
  wire n6755_o;
  wire n6757_o;
  wire n6761_o;
  wire [1:0] n6762_o;
  wire [7:0] n6763_o;
  wire [7:0] n6764_o;
  wire [7:0] n6765_o;
  wire [7:0] n6766_o;
  localparam [3:0] n6767_o = 4'b0000;
  wire [1:0] n6768_o;
  wire n6774_o;
  wire [15:0] n6775_o;
  wire [15:0] n6776_o;
  wire n6777_o;
  wire n6778_o;
  wire [3:0] n6781_o;
  wire n6783_o;
  wire [1:0] n6785_o;
  wire [7:0] n6786_o;
  wire [7:0] n6787_o;
  reg [7:0] n6788_o;
  wire [7:0] n6789_o;
  wire [7:0] n6790_o;
  reg [7:0] n6791_o;
  wire [7:0] n6792_o;
  wire [7:0] n6793_o;
  reg [7:0] n6794_o;
  wire [7:0] n6795_o;
  wire [7:0] n6796_o;
  reg [7:0] n6797_o;
  reg [3:0] n6798_o;
  wire [35:0] n6799_o;
  wire [35:0] n6804_o;
  wire n6808_o;
  wire [1:0] n6810_o;
  wire [1:0] n6811_o;
  wire [7:0] n6812_o;
  wire n6813_o;
  wire n6814_o;
  wire n6815_o;
  wire n6816_o;
  wire n6817_o;
  wire n6818_o;
  wire n6819_o;
  wire n6820_o;
  wire n6821_o;
  wire n6822_o;
  wire n6823_o;
  wire n6824_o;
  wire n6825_o;
  wire n6826_o;
  wire n6827_o;
  wire n6828_o;
  wire n6829_o;
  wire n6830_o;
  wire n6831_o;
  wire n6832_o;
  wire n6833_o;
  wire n6834_o;
  wire n6835_o;
  wire n6836_o;
  wire n6837_o;
  wire n6838_o;
  wire n6839_o;
  wire n6840_o;
  wire n6841_o;
  wire n6842_o;
  wire n6843_o;
  wire n6844_o;
  wire n6845_o;
  wire n6846_o;
  wire n6847_o;
  wire n6848_o;
  wire n6849_o;
  wire n6850_o;
  wire n6851_o;
  wire n6852_o;
  wire n6853_o;
  wire n6854_o;
  wire n6855_o;
  wire n6856_o;
  wire n6857_o;
  wire n6858_o;
  wire n6859_o;
  wire n6860_o;
  wire n6861_o;
  wire n6862_o;
  wire n6863_o;
  wire n6864_o;
  wire n6865_o;
  wire n6866_o;
  wire n6867_o;
  wire n6868_o;
  wire n6869_o;
  wire n6870_o;
  wire n6871_o;
  wire n6872_o;
  wire n6873_o;
  wire n6874_o;
  wire n6875_o;
  wire n6876_o;
  wire n6877_o;
  wire n6878_o;
  wire n6879_o;
  wire n6880_o;
  wire n6881_o;
  wire n6882_o;
  wire n6883_o;
  wire n6884_o;
  wire n6885_o;
  wire n6886_o;
  wire n6887_o;
  wire n6888_o;
  wire n6889_o;
  wire n6890_o;
  wire n6891_o;
  wire n6892_o;
  wire n6893_o;
  wire n6894_o;
  wire n6895_o;
  wire n6896_o;
  wire n6897_o;
  wire n6898_o;
  wire n6899_o;
  wire n6900_o;
  wire n6901_o;
  wire n6902_o;
  wire n6903_o;
  wire n6904_o;
  wire n6905_o;
  wire n6906_o;
  wire n6907_o;
  wire n6908_o;
  wire [3:0] n6909_o;
  wire [3:0] n6910_o;
  wire [3:0] n6911_o;
  wire [3:0] n6912_o;
  wire [3:0] n6913_o;
  wire [3:0] n6914_o;
  wire [15:0] n6915_o;
  wire [7:0] n6916_o;
  wire [23:0] n6917_o;
  wire n6919_o;
  wire [7:0] n6920_o;
  wire n6921_o;
  wire n6922_o;
  wire n6923_o;
  wire n6924_o;
  wire n6925_o;
  wire n6926_o;
  wire n6927_o;
  wire n6928_o;
  wire n6929_o;
  wire n6930_o;
  wire n6931_o;
  wire n6932_o;
  wire n6933_o;
  wire n6934_o;
  wire n6935_o;
  wire n6936_o;
  wire n6937_o;
  wire n6938_o;
  wire n6939_o;
  wire n6940_o;
  wire n6941_o;
  wire n6942_o;
  wire n6943_o;
  wire n6944_o;
  wire n6945_o;
  wire n6946_o;
  wire n6947_o;
  wire n6948_o;
  wire n6949_o;
  wire n6950_o;
  wire n6951_o;
  wire n6952_o;
  wire n6953_o;
  wire n6954_o;
  wire n6955_o;
  wire n6956_o;
  wire n6957_o;
  wire n6958_o;
  wire n6959_o;
  wire n6960_o;
  wire n6961_o;
  wire n6962_o;
  wire n6963_o;
  wire n6964_o;
  wire n6965_o;
  wire n6966_o;
  wire n6967_o;
  wire n6968_o;
  wire n6969_o;
  wire n6970_o;
  wire n6971_o;
  wire n6972_o;
  wire n6973_o;
  wire n6974_o;
  wire n6975_o;
  wire n6976_o;
  wire n6977_o;
  wire n6978_o;
  wire n6979_o;
  wire n6980_o;
  wire n6981_o;
  wire n6982_o;
  wire n6983_o;
  wire n6984_o;
  wire n6985_o;
  wire n6986_o;
  wire n6987_o;
  wire n6988_o;
  wire n6989_o;
  wire n6990_o;
  wire n6991_o;
  wire n6992_o;
  wire n6993_o;
  wire n6994_o;
  wire n6995_o;
  wire n6996_o;
  wire n6997_o;
  wire n6998_o;
  wire n6999_o;
  wire n7000_o;
  wire n7001_o;
  wire n7002_o;
  wire n7003_o;
  wire n7004_o;
  wire n7005_o;
  wire n7006_o;
  wire n7007_o;
  wire n7008_o;
  wire n7009_o;
  wire n7010_o;
  wire n7011_o;
  wire n7012_o;
  wire n7013_o;
  wire n7014_o;
  wire n7015_o;
  wire n7016_o;
  wire [3:0] n7017_o;
  wire [3:0] n7018_o;
  wire [3:0] n7019_o;
  wire [3:0] n7020_o;
  wire [3:0] n7021_o;
  wire [3:0] n7022_o;
  wire [15:0] n7023_o;
  wire [7:0] n7024_o;
  wire [23:0] n7025_o;
  wire n7027_o;
  wire [7:0] n7028_o;
  wire n7029_o;
  wire n7030_o;
  wire n7031_o;
  wire n7032_o;
  wire n7033_o;
  wire n7034_o;
  wire n7035_o;
  wire n7036_o;
  wire n7037_o;
  wire n7038_o;
  wire n7039_o;
  wire n7040_o;
  wire n7041_o;
  wire n7042_o;
  wire n7043_o;
  wire n7044_o;
  wire n7045_o;
  wire n7046_o;
  wire n7047_o;
  wire n7048_o;
  wire n7049_o;
  wire n7050_o;
  wire n7051_o;
  wire n7052_o;
  wire n7053_o;
  wire n7054_o;
  wire n7055_o;
  wire n7056_o;
  wire n7057_o;
  wire n7058_o;
  wire n7059_o;
  wire n7060_o;
  wire n7061_o;
  wire n7062_o;
  wire n7063_o;
  wire n7064_o;
  wire n7065_o;
  wire n7066_o;
  wire n7067_o;
  wire n7068_o;
  wire n7069_o;
  wire n7070_o;
  wire n7071_o;
  wire n7072_o;
  wire n7073_o;
  wire n7074_o;
  wire n7075_o;
  wire n7076_o;
  wire n7077_o;
  wire n7078_o;
  wire n7079_o;
  wire n7080_o;
  wire n7081_o;
  wire n7082_o;
  wire n7083_o;
  wire n7084_o;
  wire n7085_o;
  wire n7086_o;
  wire n7087_o;
  wire n7088_o;
  wire n7089_o;
  wire n7090_o;
  wire n7091_o;
  wire n7092_o;
  wire n7093_o;
  wire n7094_o;
  wire n7095_o;
  wire n7096_o;
  wire n7097_o;
  wire n7098_o;
  wire n7099_o;
  wire n7100_o;
  wire n7101_o;
  wire n7102_o;
  wire n7103_o;
  wire n7104_o;
  wire n7105_o;
  wire n7106_o;
  wire n7107_o;
  wire n7108_o;
  wire n7109_o;
  wire n7110_o;
  wire n7111_o;
  wire n7112_o;
  wire n7113_o;
  wire n7114_o;
  wire n7115_o;
  wire n7116_o;
  wire n7117_o;
  wire n7118_o;
  wire n7119_o;
  wire n7120_o;
  wire n7121_o;
  wire n7122_o;
  wire n7123_o;
  wire n7124_o;
  wire [3:0] n7125_o;
  wire [3:0] n7126_o;
  wire [3:0] n7127_o;
  wire [3:0] n7128_o;
  wire [3:0] n7129_o;
  wire [3:0] n7130_o;
  wire [15:0] n7131_o;
  wire [7:0] n7132_o;
  wire [23:0] n7133_o;
  wire n7135_o;
  wire [7:0] n7136_o;
  wire n7137_o;
  wire n7138_o;
  wire n7139_o;
  wire n7140_o;
  wire n7141_o;
  wire n7142_o;
  wire n7143_o;
  wire n7144_o;
  wire n7145_o;
  wire n7146_o;
  wire n7147_o;
  wire n7148_o;
  wire n7149_o;
  wire n7150_o;
  wire n7151_o;
  wire n7152_o;
  wire n7153_o;
  wire n7154_o;
  wire n7155_o;
  wire n7156_o;
  wire n7157_o;
  wire n7158_o;
  wire n7159_o;
  wire n7160_o;
  wire n7161_o;
  wire n7162_o;
  wire n7163_o;
  wire n7164_o;
  wire n7165_o;
  wire n7166_o;
  wire n7167_o;
  wire n7168_o;
  wire n7169_o;
  wire n7170_o;
  wire n7171_o;
  wire n7172_o;
  wire n7173_o;
  wire n7174_o;
  wire n7175_o;
  wire n7176_o;
  wire n7177_o;
  wire n7178_o;
  wire n7179_o;
  wire n7180_o;
  wire n7181_o;
  wire n7182_o;
  wire n7183_o;
  wire n7184_o;
  wire n7185_o;
  wire n7186_o;
  wire n7187_o;
  wire n7188_o;
  wire n7189_o;
  wire n7190_o;
  wire n7191_o;
  wire n7192_o;
  wire n7193_o;
  wire n7194_o;
  wire n7195_o;
  wire n7196_o;
  wire n7197_o;
  wire n7198_o;
  wire n7199_o;
  wire n7200_o;
  wire n7201_o;
  wire n7202_o;
  wire n7203_o;
  wire n7204_o;
  wire n7205_o;
  wire n7206_o;
  wire n7207_o;
  wire n7208_o;
  wire n7209_o;
  wire n7210_o;
  wire n7211_o;
  wire n7212_o;
  wire n7213_o;
  wire n7214_o;
  wire n7215_o;
  wire n7216_o;
  wire n7217_o;
  wire n7218_o;
  wire n7219_o;
  wire n7220_o;
  wire n7221_o;
  wire n7222_o;
  wire n7223_o;
  wire n7224_o;
  wire n7225_o;
  wire n7226_o;
  wire n7227_o;
  wire n7228_o;
  wire n7229_o;
  wire n7230_o;
  wire n7231_o;
  wire n7232_o;
  wire [3:0] n7233_o;
  wire [3:0] n7234_o;
  wire [3:0] n7235_o;
  wire [3:0] n7236_o;
  wire [3:0] n7237_o;
  wire [3:0] n7238_o;
  wire [15:0] n7239_o;
  wire [7:0] n7240_o;
  wire [23:0] n7241_o;
  wire [2:0] n7242_o;
  reg [7:0] n7243_o;
  reg [23:0] n7244_o;
  wire n7246_o;
  wire n7247_o;
  wire n7248_o;
  wire [15:0] n7249_o;
  wire n7250_o;
  wire n7251_o;
  wire n7252_o;
  wire n7253_o;
  wire n7254_o;
  wire n7255_o;
  wire n7256_o;
  wire n7257_o;
  wire n7258_o;
  wire n7259_o;
  wire n7260_o;
  wire n7261_o;
  wire n7262_o;
  wire n7263_o;
  wire n7264_o;
  wire n7265_o;
  wire n7266_o;
  wire n7267_o;
  wire n7268_o;
  wire n7269_o;
  wire n7270_o;
  wire n7271_o;
  wire n7272_o;
  wire n7273_o;
  wire n7274_o;
  wire n7275_o;
  wire n7276_o;
  wire n7277_o;
  wire n7278_o;
  wire n7279_o;
  wire n7280_o;
  wire n7281_o;
  wire n7282_o;
  wire n7283_o;
  wire n7284_o;
  wire n7285_o;
  wire n7286_o;
  wire n7287_o;
  wire n7288_o;
  wire n7289_o;
  wire n7290_o;
  wire n7291_o;
  wire n7292_o;
  wire n7293_o;
  wire n7294_o;
  wire n7295_o;
  wire n7296_o;
  wire n7297_o;
  wire n7298_o;
  wire n7299_o;
  wire n7300_o;
  wire n7301_o;
  wire n7302_o;
  wire n7303_o;
  wire n7304_o;
  wire n7305_o;
  wire n7306_o;
  wire n7307_o;
  wire n7308_o;
  wire n7309_o;
  wire n7310_o;
  wire n7311_o;
  wire n7312_o;
  wire n7313_o;
  wire [3:0] n7314_o;
  wire [3:0] n7315_o;
  wire [3:0] n7316_o;
  wire [3:0] n7317_o;
  wire [15:0] n7318_o;
  wire [15:0] n7319_o;
  wire n7320_o;
  wire n7321_o;
  wire n7322_o;
  wire n7323_o;
  wire n7324_o;
  wire n7325_o;
  wire n7326_o;
  wire n7327_o;
  wire n7328_o;
  wire n7329_o;
  wire n7330_o;
  wire n7331_o;
  wire n7332_o;
  wire n7333_o;
  wire n7334_o;
  wire n7335_o;
  wire n7336_o;
  wire n7337_o;
  wire n7338_o;
  wire n7339_o;
  wire n7340_o;
  wire n7341_o;
  wire n7342_o;
  wire n7343_o;
  wire n7344_o;
  wire n7345_o;
  wire n7346_o;
  wire n7347_o;
  wire n7348_o;
  wire n7349_o;
  wire n7350_o;
  wire n7351_o;
  wire n7352_o;
  wire n7353_o;
  wire n7354_o;
  wire n7355_o;
  wire n7356_o;
  wire n7357_o;
  wire n7358_o;
  wire n7359_o;
  wire n7360_o;
  wire n7361_o;
  wire n7362_o;
  wire n7363_o;
  wire n7364_o;
  wire n7365_o;
  wire n7366_o;
  wire n7367_o;
  wire n7368_o;
  wire n7369_o;
  wire n7370_o;
  wire n7371_o;
  wire n7372_o;
  wire n7373_o;
  wire n7374_o;
  wire n7375_o;
  wire n7376_o;
  wire n7377_o;
  wire n7378_o;
  wire n7379_o;
  wire n7380_o;
  wire n7381_o;
  wire n7382_o;
  wire n7383_o;
  wire [3:0] n7384_o;
  wire [3:0] n7385_o;
  wire [3:0] n7386_o;
  wire [3:0] n7387_o;
  wire [15:0] n7388_o;
  wire [31:0] n7389_o;
  wire [31:0] n7390_o;
  wire [31:0] n7391_o;
  wire n7393_o;
  wire [31:0] n7394_o;
  wire [1:0] n7395_o;
  wire [7:0] n7396_o;
  wire [7:0] n7397_o;
  reg [7:0] n7398_o;
  wire [23:0] n7399_o;
  wire [23:0] n7400_o;
  reg [23:0] n7401_o;
  wire [31:0] n7402_o;
  wire n7409_o;
  wire n7411_o;
  wire n7412_o;
  wire n7413_o;
  wire n7414_o;
  wire n7415_o;
  wire n7416_o;
  wire n7417_o;
  wire n7419_o;
  wire n7420_o;
  wire n7428_o;
  wire n7429_o;
  wire n7430_o;
  wire n7431_o;
  wire n7432_o;
  wire n7433_o;
  wire n7434_o;
  wire n7435_o;
  wire n7436_o;
  wire n7437_o;
  wire n7438_o;
  wire n7439_o;
  wire n7440_o;
  wire n7441_o;
  wire n7442_o;
  wire n7443_o;
  wire n7444_o;
  wire n7445_o;
  wire n7446_o;
  wire n7447_o;
  wire n7448_o;
  wire [31:0] n7449_o;
  reg [31:0] n7450_q;
  wire n7451_o;
  reg n7452_q;
  reg n7453_q;
  reg n7454_q;
  wire [31:0] n7455_o;
  reg [31:0] n7456_q;
  wire [35:0] n7457_o;
  wire [35:0] n7458_o;
  reg [35:0] n7459_q;
  wire [1:0] n7460_o;
  wire [1:0] n7461_o;
  reg [1:0] n7462_q;
  wire n7463_o;
  wire n7464_o;
  reg n7465_q;
  wire [73:0] n7466_o;
  wire n7467_o;
  wire n7468_o;
  wire n7469_o;
  wire n7470_o;
  wire n7471_o;
  wire n7472_o;
  wire n7473_o;
  wire n7474_o;
  wire n7475_o;
  wire n7476_o;
  wire n7477_o;
  wire n7478_o;
  wire n7479_o;
  wire n7480_o;
  wire n7481_o;
  wire n7482_o;
  wire [3:0] n7483_o;
  assign rdata_o = n7456_q; //(module output)
  assign mar_o = mar; //(module output)
  assign wait_o = n7429_o; //(module output)
  assign ma_load_o = n7433_o; //(module output)
  assign ma_store_o = n7440_o; //(module output)
  assign be_load_o = n7437_o; //(module output)
  assign be_store_o = n7443_o; //(module output)
  assign bus_req_o_addr = n6696_o; //(module output)
  assign bus_req_o_data = n6697_o; //(module output)
  assign bus_req_o_ben = n6698_o; //(module output)
  assign bus_req_o_stb = n6699_o; //(module output)
  assign bus_req_o_rw = n6700_o; //(module output)
  assign bus_req_o_src = n6701_o; //(module output)
  assign bus_req_o_priv = n6702_o; //(module output)
  assign bus_req_o_rvso = n6703_o; //(module output)
  assign bus_req_o_fence = n6704_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:224:18  */
  assign n6687_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_lsu_priv, ctrl_i_lsu_fence, ctrl_i_lsu_mo_we, ctrl_i_lsu_rw, ctrl_i_lsu_req, ctrl_i_alu_cp_trig, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  assign n6696_o = n7466_o[31:0]; // extract
  assign n6697_o = n7466_o[63:32]; // extract
  assign n6698_o = n7466_o[67:64]; // extract
  assign n6699_o = n7466_o[68]; // extract
  assign n6700_o = n7466_o[69]; // extract
  assign n6701_o = n7466_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:143:3  */
  assign n6702_o = n7466_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:107:22  */
  assign n6703_o = n7466_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:107:10  */
  assign n6704_o = n7466_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:106:22  */
  assign n6705_o = {bus_rsp_i_err, bus_rsp_i_ack, bus_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:69:10  */
  assign mar = n7450_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:70:10  */
  assign misaligned = n7452_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:71:10  */
  assign arbiter_req = n7453_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:72:10  */
  assign arbiter_err = n7454_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:80:16  */
  assign n6707_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:84:18  */
  assign n6709_o = n6687_o[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:86:30  */
  assign n6710_o = n6687_o[42:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:87:11  */
  assign n6712_o = n6710_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:88:46  */
  assign n6713_o = addr_i[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:88:11  */
  assign n6715_o = n6710_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:89:46  */
  assign n6716_o = addr_i[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:89:59  */
  assign n6717_o = addr_i[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:89:50  */
  assign n6718_o = n6716_o | n6717_o;
  assign n6719_o = {n6715_o, n6712_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:86:9  */
  always @*
    case (n6719_o)
      2'b10: n6721_o = n6713_o;
      2'b01: n6721_o = 1'b0;
      default: n6721_o = n6718_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:104:16  */
  assign n6732_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:109:18  */
  assign n6737_o = n6687_o[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:111:32  */
  assign n6738_o = n6687_o[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:113:34  */
  assign n6739_o = n6687_o[40]; // extract
  assign n6741_o = {1'b0, n6739_o};
  assign n6750_o = {1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:128:29  */
  assign n6755_o = n6687_o[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:135:16  */
  assign n6757_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:139:18  */
  assign n6761_o = n6687_o[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:140:30  */
  assign n6762_o = n6687_o[42:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:142:52  */
  assign n6763_o = wdata_i[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:143:52  */
  assign n6764_o = wdata_i[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:144:52  */
  assign n6765_o = wdata_i[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:145:52  */
  assign n6766_o = wdata_i[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:53  */
  assign n6768_o = addr_i[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:141:11  */
  assign n6774_o = n6762_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:149:52  */
  assign n6775_o = wdata_i[15:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:150:52  */
  assign n6776_o = wdata_i[15:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:151:23  */
  assign n6777_o = addr_i[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:151:27  */
  assign n6778_o = ~n6777_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:151:13  */
  assign n6781_o = n6778_o ? 4'b0011 : 4'b1100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:148:11  */
  assign n6783_o = n6762_o == 2'b01;
  assign n6785_o = {n6783_o, n6774_o};
  assign n6786_o = n6775_o[7:0]; // extract
  assign n6787_o = wdata_i[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:140:9  */
  always @*
    case (n6785_o)
      2'b10: n6788_o = n6786_o;
      2'b01: n6788_o = n6763_o;
      default: n6788_o = n6787_o;
    endcase
  assign n6789_o = n6775_o[15:8]; // extract
  assign n6790_o = wdata_i[15:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:140:9  */
  always @*
    case (n6785_o)
      2'b10: n6791_o = n6789_o;
      2'b01: n6791_o = n6764_o;
      default: n6791_o = n6790_o;
    endcase
  assign n6792_o = n6776_o[7:0]; // extract
  assign n6793_o = wdata_i[23:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:140:9  */
  always @*
    case (n6785_o)
      2'b10: n6794_o = n6792_o;
      2'b01: n6794_o = n6765_o;
      default: n6794_o = n6793_o;
    endcase
  assign n6795_o = n6776_o[15:8]; // extract
  assign n6796_o = wdata_i[31:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:140:9  */
  always @*
    case (n6785_o)
      2'b10: n6797_o = n6795_o;
      2'b01: n6797_o = n6766_o;
      default: n6797_o = n6796_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:140:9  */
  always @*
    case (n6785_o)
      2'b10: n6798_o = n6781_o;
      2'b01: n6798_o = n7483_o;
      default: n6798_o = 4'b1111;
    endcase
  assign n6799_o = {n6798_o, n6797_o, n6794_o, n6791_o, n6788_o};
  assign n6804_o = {4'b0000, 32'b00000000000000000000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:169:16  */
  assign n6808_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:173:30  */
  assign n6810_o = n6687_o[42:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:175:21  */
  assign n6811_o = mar[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:177:54  */
  assign n6812_o = n6705_o[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6813_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6814_o = ~n6813_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6815_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6816_o = n6814_o & n6815_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6817_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6818_o = ~n6817_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6819_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6820_o = n6818_o & n6819_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6821_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6822_o = ~n6821_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6823_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6824_o = n6822_o & n6823_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6825_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6826_o = ~n6825_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6827_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6828_o = n6826_o & n6827_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6829_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6830_o = ~n6829_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6831_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6832_o = n6830_o & n6831_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6833_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6834_o = ~n6833_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6835_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6836_o = n6834_o & n6835_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6837_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6838_o = ~n6837_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6839_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6840_o = n6838_o & n6839_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6841_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6842_o = ~n6841_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6843_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6844_o = n6842_o & n6843_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6845_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6846_o = ~n6845_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6847_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6848_o = n6846_o & n6847_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6849_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6850_o = ~n6849_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6851_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6852_o = n6850_o & n6851_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6853_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6854_o = ~n6853_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6855_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6856_o = n6854_o & n6855_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6857_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6858_o = ~n6857_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6859_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6860_o = n6858_o & n6859_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6861_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6862_o = ~n6861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6863_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6864_o = n6862_o & n6863_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6865_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6866_o = ~n6865_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6867_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6868_o = n6866_o & n6867_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6869_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6870_o = ~n6869_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6871_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6872_o = n6870_o & n6871_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6873_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6874_o = ~n6873_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6875_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6876_o = n6874_o & n6875_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6877_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6878_o = ~n6877_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6879_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6880_o = n6878_o & n6879_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6881_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6882_o = ~n6881_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6883_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6884_o = n6882_o & n6883_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6885_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6886_o = ~n6885_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6887_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6888_o = n6886_o & n6887_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6889_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6890_o = ~n6889_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6891_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6892_o = n6890_o & n6891_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6893_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6894_o = ~n6893_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6895_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6896_o = n6894_o & n6895_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6897_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6898_o = ~n6897_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6899_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6900_o = n6898_o & n6899_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6901_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6902_o = ~n6901_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6903_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6904_o = n6902_o & n6903_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:78  */
  assign n6905_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:58  */
  assign n6906_o = ~n6905_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:101  */
  assign n6907_o = n6705_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:178:83  */
  assign n6908_o = n6906_o & n6907_o;
  assign n6909_o = {n6816_o, n6820_o, n6824_o, n6828_o};
  assign n6910_o = {n6832_o, n6836_o, n6840_o, n6844_o};
  assign n6911_o = {n6848_o, n6852_o, n6856_o, n6860_o};
  assign n6912_o = {n6864_o, n6868_o, n6872_o, n6876_o};
  assign n6913_o = {n6880_o, n6884_o, n6888_o, n6892_o};
  assign n6914_o = {n6896_o, n6900_o, n6904_o, n6908_o};
  assign n6915_o = {n6909_o, n6910_o, n6911_o, n6912_o};
  assign n6916_o = {n6913_o, n6914_o};
  assign n6917_o = {n6915_o, n6916_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:176:15  */
  assign n6919_o = n6811_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:180:54  */
  assign n6920_o = n6705_o[15:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6921_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6922_o = ~n6921_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6923_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6924_o = n6922_o & n6923_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6925_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6926_o = ~n6925_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6927_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6928_o = n6926_o & n6927_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6929_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6930_o = ~n6929_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6931_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6932_o = n6930_o & n6931_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6933_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6934_o = ~n6933_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6935_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6936_o = n6934_o & n6935_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6937_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6938_o = ~n6937_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6939_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6940_o = n6938_o & n6939_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6941_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6942_o = ~n6941_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6943_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6944_o = n6942_o & n6943_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6945_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6946_o = ~n6945_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6947_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6948_o = n6946_o & n6947_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6949_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6950_o = ~n6949_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6951_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6952_o = n6950_o & n6951_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6953_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6954_o = ~n6953_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6955_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6956_o = n6954_o & n6955_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6957_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6958_o = ~n6957_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6959_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6960_o = n6958_o & n6959_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6961_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6962_o = ~n6961_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6963_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6964_o = n6962_o & n6963_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6965_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6966_o = ~n6965_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6967_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6968_o = n6966_o & n6967_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6969_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6970_o = ~n6969_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6971_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6972_o = n6970_o & n6971_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6973_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6974_o = ~n6973_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6975_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6976_o = n6974_o & n6975_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6977_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6978_o = ~n6977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6979_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6980_o = n6978_o & n6979_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6981_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6982_o = ~n6981_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6983_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6984_o = n6982_o & n6983_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6985_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6986_o = ~n6985_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6987_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6988_o = n6986_o & n6987_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6989_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6990_o = ~n6989_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6991_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6992_o = n6990_o & n6991_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6993_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6994_o = ~n6993_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6995_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n6996_o = n6994_o & n6995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n6997_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n6998_o = ~n6997_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n6999_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n7000_o = n6998_o & n6999_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n7001_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n7002_o = ~n7001_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n7003_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n7004_o = n7002_o & n7003_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n7005_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n7006_o = ~n7005_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n7007_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n7008_o = n7006_o & n7007_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n7009_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n7010_o = ~n7009_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n7011_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n7012_o = n7010_o & n7011_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:78  */
  assign n7013_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:58  */
  assign n7014_o = ~n7013_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:101  */
  assign n7015_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:181:83  */
  assign n7016_o = n7014_o & n7015_o;
  assign n7017_o = {n6924_o, n6928_o, n6932_o, n6936_o};
  assign n7018_o = {n6940_o, n6944_o, n6948_o, n6952_o};
  assign n7019_o = {n6956_o, n6960_o, n6964_o, n6968_o};
  assign n7020_o = {n6972_o, n6976_o, n6980_o, n6984_o};
  assign n7021_o = {n6988_o, n6992_o, n6996_o, n7000_o};
  assign n7022_o = {n7004_o, n7008_o, n7012_o, n7016_o};
  assign n7023_o = {n7017_o, n7018_o, n7019_o, n7020_o};
  assign n7024_o = {n7021_o, n7022_o};
  assign n7025_o = {n7023_o, n7024_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:179:15  */
  assign n7027_o = n6811_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:183:54  */
  assign n7028_o = n6705_o[23:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7029_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7030_o = ~n7029_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7031_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7032_o = n7030_o & n7031_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7033_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7034_o = ~n7033_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7035_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7036_o = n7034_o & n7035_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7037_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7038_o = ~n7037_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7039_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7040_o = n7038_o & n7039_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7041_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7042_o = ~n7041_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7043_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7044_o = n7042_o & n7043_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7045_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7046_o = ~n7045_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7047_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7048_o = n7046_o & n7047_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7049_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7050_o = ~n7049_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7051_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7052_o = n7050_o & n7051_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7053_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7054_o = ~n7053_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7055_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7056_o = n7054_o & n7055_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7057_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7058_o = ~n7057_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7059_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7060_o = n7058_o & n7059_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7061_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7062_o = ~n7061_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7063_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7064_o = n7062_o & n7063_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7065_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7066_o = ~n7065_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7067_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7068_o = n7066_o & n7067_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7069_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7070_o = ~n7069_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7071_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7072_o = n7070_o & n7071_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7073_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7074_o = ~n7073_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7075_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7076_o = n7074_o & n7075_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7077_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7078_o = ~n7077_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7079_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7080_o = n7078_o & n7079_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7081_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7082_o = ~n7081_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7083_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7084_o = n7082_o & n7083_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7085_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7086_o = ~n7085_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7087_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7088_o = n7086_o & n7087_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7089_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7090_o = ~n7089_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7091_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7092_o = n7090_o & n7091_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7093_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7094_o = ~n7093_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7095_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7096_o = n7094_o & n7095_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7097_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7098_o = ~n7097_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7099_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7100_o = n7098_o & n7099_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7101_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7102_o = ~n7101_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7103_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7104_o = n7102_o & n7103_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7105_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7106_o = ~n7105_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7107_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7108_o = n7106_o & n7107_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7109_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7110_o = ~n7109_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7111_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7112_o = n7110_o & n7111_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7113_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7114_o = ~n7113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7115_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7116_o = n7114_o & n7115_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7117_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7118_o = ~n7117_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7119_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7120_o = n7118_o & n7119_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:78  */
  assign n7121_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:58  */
  assign n7122_o = ~n7121_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:101  */
  assign n7123_o = n6705_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:184:83  */
  assign n7124_o = n7122_o & n7123_o;
  assign n7125_o = {n7032_o, n7036_o, n7040_o, n7044_o};
  assign n7126_o = {n7048_o, n7052_o, n7056_o, n7060_o};
  assign n7127_o = {n7064_o, n7068_o, n7072_o, n7076_o};
  assign n7128_o = {n7080_o, n7084_o, n7088_o, n7092_o};
  assign n7129_o = {n7096_o, n7100_o, n7104_o, n7108_o};
  assign n7130_o = {n7112_o, n7116_o, n7120_o, n7124_o};
  assign n7131_o = {n7125_o, n7126_o, n7127_o, n7128_o};
  assign n7132_o = {n7129_o, n7130_o};
  assign n7133_o = {n7131_o, n7132_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:182:15  */
  assign n7135_o = n6811_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:186:54  */
  assign n7136_o = n6705_o[31:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7137_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7138_o = ~n7137_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7139_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7140_o = n7138_o & n7139_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7141_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7142_o = ~n7141_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7143_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7144_o = n7142_o & n7143_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7145_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7146_o = ~n7145_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7147_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7148_o = n7146_o & n7147_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7149_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7150_o = ~n7149_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7151_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7152_o = n7150_o & n7151_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7153_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7154_o = ~n7153_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7155_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7156_o = n7154_o & n7155_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7157_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7158_o = ~n7157_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7159_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7160_o = n7158_o & n7159_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7161_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7162_o = ~n7161_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7163_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7164_o = n7162_o & n7163_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7165_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7166_o = ~n7165_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7167_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7168_o = n7166_o & n7167_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7169_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7170_o = ~n7169_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7171_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7172_o = n7170_o & n7171_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7173_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7174_o = ~n7173_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7175_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7176_o = n7174_o & n7175_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7177_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7178_o = ~n7177_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7179_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7180_o = n7178_o & n7179_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7181_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7182_o = ~n7181_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7183_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7184_o = n7182_o & n7183_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7185_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7186_o = ~n7185_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7187_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7188_o = n7186_o & n7187_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7189_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7190_o = ~n7189_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7191_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7192_o = n7190_o & n7191_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7193_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7194_o = ~n7193_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7195_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7196_o = n7194_o & n7195_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7197_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7198_o = ~n7197_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7199_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7200_o = n7198_o & n7199_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7201_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7202_o = ~n7201_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7203_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7204_o = n7202_o & n7203_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7205_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7206_o = ~n7205_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7207_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7208_o = n7206_o & n7207_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7209_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7210_o = ~n7209_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7211_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7212_o = n7210_o & n7211_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7213_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7214_o = ~n7213_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7215_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7216_o = n7214_o & n7215_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7217_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7218_o = ~n7217_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7219_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7220_o = n7218_o & n7219_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7221_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7222_o = ~n7221_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7223_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7224_o = n7222_o & n7223_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7225_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7226_o = ~n7225_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7227_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7228_o = n7226_o & n7227_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:78  */
  assign n7229_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:58  */
  assign n7230_o = ~n7229_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:101  */
  assign n7231_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:187:83  */
  assign n7232_o = n7230_o & n7231_o;
  assign n7233_o = {n7140_o, n7144_o, n7148_o, n7152_o};
  assign n7234_o = {n7156_o, n7160_o, n7164_o, n7168_o};
  assign n7235_o = {n7172_o, n7176_o, n7180_o, n7184_o};
  assign n7236_o = {n7188_o, n7192_o, n7196_o, n7200_o};
  assign n7237_o = {n7204_o, n7208_o, n7212_o, n7216_o};
  assign n7238_o = {n7220_o, n7224_o, n7228_o, n7232_o};
  assign n7239_o = {n7233_o, n7234_o, n7235_o, n7236_o};
  assign n7240_o = {n7237_o, n7238_o};
  assign n7241_o = {n7239_o, n7240_o};
  assign n7242_o = {n7135_o, n7027_o, n6919_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:175:13  */
  always @*
    case (n7242_o)
      3'b100: n7243_o = n7028_o;
      3'b010: n7243_o = n6920_o;
      3'b001: n7243_o = n6812_o;
      default: n7243_o = n7136_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:175:13  */
  always @*
    case (n7242_o)
      3'b100: n7244_o = n7133_o;
      3'b010: n7244_o = n7025_o;
      3'b001: n7244_o = n6917_o;
      default: n7244_o = n7241_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:174:11  */
  assign n7246_o = n6810_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:190:20  */
  assign n7247_o = mar[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:190:24  */
  assign n7248_o = ~n7247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:191:53  */
  assign n7249_o = n6705_o[15:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7250_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7251_o = ~n7250_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7252_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7253_o = n7251_o & n7252_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7254_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7255_o = ~n7254_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7256_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7257_o = n7255_o & n7256_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7258_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7259_o = ~n7258_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7260_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7261_o = n7259_o & n7260_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7262_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7263_o = ~n7262_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7264_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7265_o = n7263_o & n7264_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7266_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7267_o = ~n7266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7268_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7269_o = n7267_o & n7268_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7270_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7271_o = ~n7270_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7272_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7273_o = n7271_o & n7272_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7274_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7275_o = ~n7274_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7276_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7277_o = n7275_o & n7276_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7278_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7279_o = ~n7278_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7280_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7281_o = n7279_o & n7280_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7282_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7283_o = ~n7282_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7284_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7285_o = n7283_o & n7284_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7286_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7287_o = ~n7286_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7288_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7289_o = n7287_o & n7288_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7290_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7291_o = ~n7290_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7292_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7293_o = n7291_o & n7292_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7294_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7295_o = ~n7294_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7296_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7297_o = n7295_o & n7296_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7298_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7299_o = ~n7298_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7300_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7301_o = n7299_o & n7300_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7302_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7303_o = ~n7302_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7304_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7305_o = n7303_o & n7304_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7306_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7307_o = ~n7306_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7308_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7309_o = n7307_o & n7308_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:77  */
  assign n7310_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:57  */
  assign n7311_o = ~n7310_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:100  */
  assign n7312_o = n6705_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:192:82  */
  assign n7313_o = n7311_o & n7312_o;
  assign n7314_o = {n7253_o, n7257_o, n7261_o, n7265_o};
  assign n7315_o = {n7269_o, n7273_o, n7277_o, n7281_o};
  assign n7316_o = {n7285_o, n7289_o, n7293_o, n7297_o};
  assign n7317_o = {n7301_o, n7305_o, n7309_o, n7313_o};
  assign n7318_o = {n7314_o, n7315_o, n7316_o, n7317_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:194:53  */
  assign n7319_o = n6705_o[31:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7320_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7321_o = ~n7320_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7322_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7323_o = n7321_o & n7322_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7324_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7325_o = ~n7324_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7326_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7327_o = n7325_o & n7326_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7328_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7329_o = ~n7328_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7330_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7331_o = n7329_o & n7330_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7332_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7333_o = ~n7332_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7334_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7335_o = n7333_o & n7334_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7336_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7337_o = ~n7336_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7338_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7339_o = n7337_o & n7338_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7340_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7341_o = ~n7340_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7342_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7343_o = n7341_o & n7342_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7344_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7345_o = ~n7344_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7346_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7347_o = n7345_o & n7346_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7348_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7349_o = ~n7348_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7350_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7351_o = n7349_o & n7350_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7352_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7353_o = ~n7352_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7354_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7355_o = n7353_o & n7354_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7356_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7357_o = ~n7356_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7358_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7359_o = n7357_o & n7358_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7360_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7361_o = ~n7360_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7362_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7363_o = n7361_o & n7362_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7364_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7365_o = ~n7364_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7366_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7367_o = n7365_o & n7366_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7368_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7369_o = ~n7368_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7370_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7371_o = n7369_o & n7370_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7372_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7373_o = ~n7372_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7374_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7375_o = n7373_o & n7374_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7376_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7377_o = ~n7376_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7378_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7379_o = n7377_o & n7378_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:77  */
  assign n7380_o = n6687_o[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:57  */
  assign n7381_o = ~n7380_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:100  */
  assign n7382_o = n6705_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:195:82  */
  assign n7383_o = n7381_o & n7382_o;
  assign n7384_o = {n7323_o, n7327_o, n7331_o, n7335_o};
  assign n7385_o = {n7339_o, n7343_o, n7347_o, n7351_o};
  assign n7386_o = {n7355_o, n7359_o, n7363_o, n7367_o};
  assign n7387_o = {n7371_o, n7375_o, n7379_o, n7383_o};
  assign n7388_o = {n7384_o, n7385_o, n7386_o, n7387_o};
  assign n7389_o = {n7388_o, n7319_o};
  assign n7390_o = {n7318_o, n7249_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:190:13  */
  assign n7391_o = n7248_o ? n7390_o : n7389_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:189:11  */
  assign n7393_o = n6810_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:198:55  */
  assign n7394_o = n6705_o[31:0]; // extract
  assign n7395_o = {n7393_o, n7246_o};
  assign n7396_o = n7391_o[7:0]; // extract
  assign n7397_o = n7394_o[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:173:9  */
  always @*
    case (n7395_o)
      2'b10: n7398_o = n7396_o;
      2'b01: n7398_o = n7243_o;
      default: n7398_o = n7397_o;
    endcase
  assign n7399_o = n7391_o[31:8]; // extract
  assign n7400_o = n7394_o[31:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:173:9  */
  always @*
    case (n7395_o)
      2'b10: n7401_o = n7399_o;
      2'b01: n7401_o = n7244_o;
      default: n7401_o = n7400_o;
    endcase
  assign n7402_o = {n7401_o, n7398_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:209:16  */
  assign n7409_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:213:32  */
  assign n7411_o = n6705_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:213:36  */
  assign n7412_o = n7411_o | pmp_fault_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:214:23  */
  assign n7413_o = ~arbiter_req;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:215:31  */
  assign n7414_o = n6687_o[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:216:24  */
  assign n7415_o = n6705_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:216:46  */
  assign n7416_o = n6687_o[65]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:216:35  */
  assign n7417_o = n7415_o | n7416_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:216:7  */
  assign n7419_o = n7417_o ? 1'b0 : arbiter_req;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:214:7  */
  assign n7420_o = n7413_o ? n7414_o : n7419_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:223:27  */
  assign n7428_o = n6705_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:223:13  */
  assign n7429_o = ~n7428_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:226:45  */
  assign n7430_o = n6687_o[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:226:34  */
  assign n7431_o = ~n7430_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:226:29  */
  assign n7432_o = arbiter_req & n7431_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:226:53  */
  assign n7433_o = n7432_o & misaligned;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:227:45  */
  assign n7434_o = n6687_o[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:227:34  */
  assign n7435_o = ~n7434_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:227:29  */
  assign n7436_o = arbiter_req & n7435_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:227:53  */
  assign n7437_o = n7436_o & arbiter_err;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:228:45  */
  assign n7438_o = n6687_o[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:228:29  */
  assign n7439_o = arbiter_req & n7438_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:228:53  */
  assign n7440_o = n7439_o & misaligned;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:229:45  */
  assign n7441_o = n6687_o[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:229:29  */
  assign n7442_o = arbiter_req & n7441_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:229:53  */
  assign n7443_o = n7442_o & arbiter_err;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:232:27  */
  assign n7444_o = n6687_o[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:232:40  */
  assign n7445_o = ~misaligned;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:232:35  */
  assign n7446_o = n7444_o & n7445_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:232:61  */
  assign n7447_o = ~pmp_fault_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:232:56  */
  assign n7448_o = n7446_o & n7447_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:83:5  */
  assign n7449_o = n6709_o ? addr_i : mar;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:83:5  */
  always @(posedge clk_i or posedge n6707_o)
    if (n6707_o)
      n7450_q <= 32'b00000000000000000000000000000000;
    else
      n7450_q <= n7449_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:83:5  */
  assign n7451_o = n6709_o ? n6721_o : misaligned;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:83:5  */
  always @(posedge clk_i or posedge n6707_o)
    if (n6707_o)
      n7452_q <= 1'b0;
    else
      n7452_q <= n7451_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:212:5  */
  always @(posedge clk_i or posedge n7409_o)
    if (n7409_o)
      n7453_q <= 1'b0;
    else
      n7453_q <= n7420_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:212:5  */
  always @(posedge clk_i or posedge n7409_o)
    if (n7409_o)
      n7454_q <= 1'b0;
    else
      n7454_q <= n7412_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:171:5  */
  assign n7455_o = arbiter_req ? n7402_o : n7456_q;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:171:5  */
  always @(posedge clk_i or posedge n6808_o)
    if (n6808_o)
      n7456_q <= 32'b00000000000000000000000000000000;
    else
      n7456_q <= n7455_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:138:5  */
  assign n7457_o = n7466_o[67:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:138:5  */
  assign n7458_o = n6761_o ? n6799_o : n7457_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:138:5  */
  always @(posedge clk_i or posedge n6757_o)
    if (n6757_o)
      n7459_q <= n6804_o;
    else
      n7459_q <= n7458_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:108:5  */
  assign n7460_o = n7466_o[72:71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:108:5  */
  assign n7461_o = n6737_o ? n6741_o : n7460_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:108:5  */
  always @(posedge clk_i or posedge n6732_o)
    if (n6732_o)
      n7462_q <= n6750_o;
    else
      n7462_q <= n7461_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:108:5  */
  assign n7463_o = n7466_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:108:5  */
  assign n7464_o = n6737_o ? n6738_o : n7463_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:108:5  */
  always @(posedge clk_i or posedge n6732_o)
    if (n6732_o)
      n7465_q <= 1'b0;
    else
      n7465_q <= n7464_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:104:5  */
  assign n7466_o = {n6755_o, n7462_q, 1'b0, n7465_q, n7448_o, n7459_q, mar};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7467_o = n6768_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7468_o = ~n7467_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7469_o = n6768_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7470_o = ~n7469_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7471_o = n7468_o & n7470_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7472_o = n7468_o & n7469_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7473_o = n7467_o & n7470_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7474_o = n7467_o & n7469_o;
  assign n7475_o = n6767_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7476_o = n7471_o ? 1'b1 : n7475_o;
  assign n7477_o = n6767_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7478_o = n7472_o ? 1'b1 : n7477_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:167:3  */
  assign n7479_o = n6767_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7480_o = n7473_o ? 1'b1 : n7479_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:138:5  */
  assign n7481_o = n6767_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_lsu.vhd:147:13  */
  assign n7482_o = n7474_o ? 1'b1 : n7481_o;
  assign n7483_o = {n7482_o, n7480_o, n7478_o, n7476_o};
endmodule

module neorv32_cpu_alu_1db721083c34eba714927c673b29edb8e81e05fb
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_lsu_req,
   input  ctrl_i_lsu_rw,
   input  ctrl_i_lsu_mo_we,
   input  ctrl_i_lsu_fence,
   input  ctrl_i_lsu_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  csr_we_i,
   input  [11:0] csr_addr_i,
   input  [31:0] csr_wdata_i,
   input  [31:0] rs1_i,
   input  [31:0] rs2_i,
   input  [31:0] rs3_i,
   input  [31:0] rs4_i,
   input  [31:0] pc_i,
   input  [31:0] imm_i,
   output [31:0] csr_rdata_o,
   output [1:0] cmp_o,
   output [31:0] res_o,
   output [31:0] add_o,
   output cp_done_o);
  wire [66:0] n6498_o;
  wire [32:0] cmp_rs1;
  wire [32:0] cmp_rs2;
  wire [1:0] cmp;
  wire [31:0] opa;
  wire [31:0] opb;
  wire [32:0] opa_x;
  wire [32:0] opb_x;
  wire [32:0] addsub_res;
  wire [31:0] cp_res;
  wire [191:0] cp_result;
  wire [5:0] cp_start;
  wire [5:0] cp_valid;
  wire [4:0] cp_shamt;
  wire [31:0] csr_rdata_fpu;
  wire [31:0] csr_rdata_cfu;
  wire n6504_o;
  wire n6505_o;
  wire n6506_o;
  wire n6507_o;
  wire [32:0] n6508_o;
  wire n6509_o;
  wire n6510_o;
  wire n6511_o;
  wire n6512_o;
  wire [32:0] n6513_o;
  wire n6515_o;
  wire n6516_o;
  wire n6519_o;
  wire n6520_o;
  wire n6522_o;
  wire [31:0] n6523_o;
  wire n6524_o;
  wire [31:0] n6525_o;
  wire n6526_o;
  wire n6527_o;
  wire n6528_o;
  wire n6529_o;
  wire [32:0] n6530_o;
  wire n6531_o;
  wire n6532_o;
  wire n6533_o;
  wire n6534_o;
  wire [32:0] n6535_o;
  wire [32:0] n6536_o;
  wire n6537_o;
  wire [32:0] n6538_o;
  wire [32:0] n6539_o;
  wire [31:0] n6540_o;
  wire [2:0] n6542_o;
  wire [31:0] n6543_o;
  wire n6545_o;
  wire [31:0] n6546_o;
  wire n6548_o;
  wire n6550_o;
  wire n6552_o;
  wire n6554_o;
  wire n6556_o;
  wire [31:0] n6557_o;
  wire n6559_o;
  wire [31:0] n6560_o;
  wire n6562_o;
  wire [31:0] n6563_o;
  wire n6565_o;
  wire [31:0] n6566_o;
  wire [7:0] n6567_o;
  wire n6568_o;
  wire n6569_o;
  wire n6570_o;
  wire n6571_o;
  wire n6572_o;
  wire n6573_o;
  wire n6574_o;
  wire n6575_o;
  reg n6576_o;
  wire [30:0] n6577_o;
  wire [30:0] n6578_o;
  wire [30:0] n6579_o;
  wire [30:0] n6580_o;
  wire [30:0] n6581_o;
  wire [30:0] n6582_o;
  wire [30:0] n6583_o;
  wire [30:0] n6584_o;
  reg [30:0] n6585_o;
  wire [5:0] n6587_o;
  wire n6588_o;
  wire n6589_o;
  wire n6590_o;
  wire n6591_o;
  wire n6592_o;
  wire n6593_o;
  wire n6594_o;
  wire n6595_o;
  wire n6596_o;
  wire n6597_o;
  wire n6598_o;
  wire [31:0] n6599_o;
  wire [31:0] n6600_o;
  wire [31:0] n6601_o;
  wire [31:0] n6602_o;
  wire [31:0] n6603_o;
  wire [31:0] n6604_o;
  wire [31:0] n6605_o;
  wire [31:0] n6606_o;
  wire [31:0] n6607_o;
  wire [31:0] n6608_o;
  wire [31:0] n6609_o;
  wire [31:0] n6610_o;
  wire [4:0] n6612_o;
  wire [31:0] neorv32_cpu_cp_shifter_inst_res_o;
  wire neorv32_cpu_cp_shifter_inst_valid_o;
  wire n6613_o;
  wire [4:0] n6614_o;
  wire [4:0] n6615_o;
  wire [4:0] n6616_o;
  wire [4:0] n6617_o;
  wire [1:0] n6618_o;
  wire n6619_o;
  wire [2:0] n6620_o;
  wire n6621_o;
  wire n6622_o;
  wire n6623_o;
  wire [5:0] n6624_o;
  wire n6625_o;
  wire n6626_o;
  wire n6627_o;
  wire n6628_o;
  wire n6629_o;
  wire [2:0] n6630_o;
  wire [11:0] n6631_o;
  wire [6:0] n6632_o;
  wire n6633_o;
  wire n6634_o;
  wire n6635_o;
  wire n6636_o;
  wire n6637_o;
  wire [31:0] neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_res_o;
  wire neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_valid_o;
  wire n6640_o;
  wire [4:0] n6641_o;
  wire [4:0] n6642_o;
  wire [4:0] n6643_o;
  wire [4:0] n6644_o;
  wire [1:0] n6645_o;
  wire n6646_o;
  wire [2:0] n6647_o;
  wire n6648_o;
  wire n6649_o;
  wire n6650_o;
  wire [5:0] n6651_o;
  wire n6652_o;
  wire n6653_o;
  wire n6654_o;
  wire n6655_o;
  wire n6656_o;
  wire [2:0] n6657_o;
  wire [11:0] n6658_o;
  wire [6:0] n6659_o;
  wire n6660_o;
  wire n6661_o;
  wire n6662_o;
  wire n6663_o;
  wire n6664_o;
  wire [1:0] n6677_o;
  wire [191:0] n6678_o;
  wire [5:0] n6679_o;
  wire [31:0] n6686_o;
  assign csr_rdata_o = n6610_o; //(module output)
  assign cmp_o = cmp; //(module output)
  assign res_o = n6686_o; //(module output)
  assign add_o = n6540_o; //(module output)
  assign cp_done_o = n6598_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:126:7  */
  assign n6498_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_lsu_priv, ctrl_i_lsu_fence, ctrl_i_lsu_mo_we, ctrl_i_lsu_rw, ctrl_i_lsu_req, ctrl_i_alu_cp_trig, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:85:10  */
  assign cmp_rs1 = n6508_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:86:10  */
  assign cmp_rs2 = n6513_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:87:10  */
  assign cmp = n6677_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:90:10  */
  assign opa = n6523_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:90:17  */
  assign opb = n6525_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:91:10  */
  assign opa_x = n6530_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:91:17  */
  assign opb_x = n6535_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:94:10  */
  assign addsub_res = n6538_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:95:10  */
  assign cp_res = n6609_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:99:10  */
  assign cp_result = n6678_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:100:10  */
  assign cp_start = n6587_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:101:10  */
  assign cp_valid = n6679_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:102:10  */
  assign cp_shamt = n6612_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:110:10  */
  assign csr_rdata_fpu = 32'b00000000000000000000000000000000; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:110:25  */
  assign csr_rdata_cfu = 32'b00000000000000000000000000000000; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:116:20  */
  assign n6504_o = rs1_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:116:49  */
  assign n6505_o = n6498_o[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:116:38  */
  assign n6506_o = ~n6505_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:116:33  */
  assign n6507_o = n6504_o & n6506_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:116:64  */
  assign n6508_o = {n6507_o, rs1_i};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:117:20  */
  assign n6509_o = rs2_i[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:117:49  */
  assign n6510_o = n6498_o[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:117:38  */
  assign n6511_o = ~n6510_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:117:33  */
  assign n6512_o = n6509_o & n6511_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:117:64  */
  assign n6513_o = {n6512_o, rs2_i};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:119:39  */
  assign n6515_o = rs1_i == rs2_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:119:27  */
  assign n6516_o = n6515_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:120:49  */
  assign n6519_o = $signed(cmp_rs1) < $signed(cmp_rs2);
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:120:27  */
  assign n6520_o = n6519_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:126:29  */
  assign n6522_o = n6498_o[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:126:16  */
  assign n6523_o = n6522_o ? pc_i : rs1_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:127:29  */
  assign n6524_o = n6498_o[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:127:16  */
  assign n6525_o = n6524_o ? imm_i : rs2_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:132:16  */
  assign n6526_o = opa[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:132:43  */
  assign n6527_o = n6498_o[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:132:32  */
  assign n6528_o = ~n6527_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:132:27  */
  assign n6529_o = n6526_o & n6528_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:132:58  */
  assign n6530_o = {n6529_o, opa};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:133:16  */
  assign n6531_o = opb[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:133:43  */
  assign n6532_o = n6498_o[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:133:32  */
  assign n6533_o = ~n6532_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:133:27  */
  assign n6534_o = n6531_o & n6533_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:133:58  */
  assign n6535_o = {n6534_o, opb};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:135:51  */
  assign n6536_o = opa_x - opb_x;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:135:89  */
  assign n6537_o = n6498_o[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:135:70  */
  assign n6538_o = n6537_o ? n6536_o : n6539_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:136:51  */
  assign n6539_o = opa_x + opb_x;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:138:22  */
  assign n6540_o = addsub_res[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:145:17  */
  assign n6542_o = n6498_o[26:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:146:48  */
  assign n6543_o = addsub_res[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:146:7  */
  assign n6545_o = n6542_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:147:48  */
  assign n6546_o = addsub_res[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:147:7  */
  assign n6548_o = n6542_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:148:7  */
  assign n6550_o = n6542_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:150:51  */
  assign n6552_o = addsub_res[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:149:7  */
  assign n6554_o = n6542_o == 3'b011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:151:7  */
  assign n6556_o = n6542_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:152:42  */
  assign n6557_o = opb ^ rs1_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:152:7  */
  assign n6559_o = n6542_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:153:42  */
  assign n6560_o = opb | rs1_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:153:7  */
  assign n6562_o = n6542_o == 3'b110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:154:42  */
  assign n6563_o = opb & rs1_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:154:7  */
  assign n6565_o = n6542_o == 3'b111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:155:48  */
  assign n6566_o = addsub_res[31:0]; // extract
  assign n6567_o = {n6565_o, n6562_o, n6559_o, n6556_o, n6554_o, n6550_o, n6548_o, n6545_o};
  assign n6568_o = n6543_o[0]; // extract
  assign n6569_o = n6546_o[0]; // extract
  assign n6570_o = cp_res[0]; // extract
  assign n6571_o = opb[0]; // extract
  assign n6572_o = n6557_o[0]; // extract
  assign n6573_o = n6560_o[0]; // extract
  assign n6574_o = n6563_o[0]; // extract
  assign n6575_o = n6566_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:145:5  */
  always @*
    case (n6567_o)
      8'b10000000: n6576_o = n6574_o;
      8'b01000000: n6576_o = n6573_o;
      8'b00100000: n6576_o = n6572_o;
      8'b00010000: n6576_o = n6571_o;
      8'b00001000: n6576_o = n6552_o;
      8'b00000100: n6576_o = n6570_o;
      8'b00000010: n6576_o = n6569_o;
      8'b00000001: n6576_o = n6568_o;
      default: n6576_o = n6575_o;
    endcase
  assign n6577_o = n6543_o[31:1]; // extract
  assign n6578_o = n6546_o[31:1]; // extract
  assign n6579_o = cp_res[31:1]; // extract
  assign n6580_o = opb[31:1]; // extract
  assign n6581_o = n6557_o[31:1]; // extract
  assign n6582_o = n6560_o[31:1]; // extract
  assign n6583_o = n6563_o[31:1]; // extract
  assign n6584_o = n6566_o[31:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:145:5  */
  always @*
    case (n6567_o)
      8'b10000000: n6585_o = n6583_o;
      8'b01000000: n6585_o = n6582_o;
      8'b00100000: n6585_o = n6581_o;
      8'b00010000: n6585_o = n6580_o;
      8'b00001000: n6585_o = 31'b0000000000000000000000000000000;
      8'b00000100: n6585_o = n6579_o;
      8'b00000010: n6585_o = n6578_o;
      8'b00000001: n6585_o = n6577_o;
      default: n6585_o = n6584_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:166:22  */
  assign n6587_o = n6498_o[35:30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:24  */
  assign n6588_o = cp_valid[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:39  */
  assign n6589_o = cp_valid[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:28  */
  assign n6590_o = n6588_o | n6589_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:54  */
  assign n6591_o = cp_valid[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:43  */
  assign n6592_o = n6590_o | n6591_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:69  */
  assign n6593_o = cp_valid[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:58  */
  assign n6594_o = n6592_o | n6593_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:84  */
  assign n6595_o = cp_valid[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:73  */
  assign n6596_o = n6594_o | n6595_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:99  */
  assign n6597_o = cp_valid[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:170:88  */
  assign n6598_o = n6596_o | n6597_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:22  */
  assign n6599_o = cp_result[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:38  */
  assign n6600_o = cp_result[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:26  */
  assign n6601_o = n6599_o | n6600_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:54  */
  assign n6602_o = cp_result[95:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:42  */
  assign n6603_o = n6601_o | n6602_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:70  */
  assign n6604_o = cp_result[127:96]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:58  */
  assign n6605_o = n6603_o | n6604_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:86  */
  assign n6606_o = cp_result[159:128]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:74  */
  assign n6607_o = n6605_o | n6606_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:102  */
  assign n6608_o = cp_result[191:160]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:174:90  */
  assign n6609_o = n6607_o | n6608_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:178:32  */
  assign n6610_o = csr_rdata_fpu | csr_rdata_cfu;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:181:18  */
  assign n6612_o = opb[4:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:186:3  */
  neorv32_cpu_cp_shifter_bf8b4530d8d246dd74ac53a13471bba17941dff7 neorv32_cpu_cp_shifter_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n6613_o),
    .ctrl_i_rf_rs1(n6614_o),
    .ctrl_i_rf_rs2(n6615_o),
    .ctrl_i_rf_rs3(n6616_o),
    .ctrl_i_rf_rd(n6617_o),
    .ctrl_i_rf_mux(n6618_o),
    .ctrl_i_rf_zero_we(n6619_o),
    .ctrl_i_alu_op(n6620_o),
    .ctrl_i_alu_opa_mux(n6621_o),
    .ctrl_i_alu_opb_mux(n6622_o),
    .ctrl_i_alu_unsigned(n6623_o),
    .ctrl_i_alu_cp_trig(n6624_o),
    .ctrl_i_lsu_req(n6625_o),
    .ctrl_i_lsu_rw(n6626_o),
    .ctrl_i_lsu_mo_we(n6627_o),
    .ctrl_i_lsu_fence(n6628_o),
    .ctrl_i_lsu_priv(n6629_o),
    .ctrl_i_ir_funct3(n6630_o),
    .ctrl_i_ir_funct12(n6631_o),
    .ctrl_i_ir_opcode(n6632_o),
    .ctrl_i_cpu_priv(n6633_o),
    .ctrl_i_cpu_sleep(n6634_o),
    .ctrl_i_cpu_trap(n6635_o),
    .ctrl_i_cpu_debug(n6636_o),
    .start_i(n6637_o),
    .rs1_i(rs1_i),
    .shamt_i(cp_shamt),
    .res_o(neorv32_cpu_cp_shifter_inst_res_o),
    .valid_o(neorv32_cpu_cp_shifter_inst_valid_o));
  assign n6613_o = n6498_o[0]; // extract
  assign n6614_o = n6498_o[5:1]; // extract
  assign n6615_o = n6498_o[10:6]; // extract
  assign n6616_o = n6498_o[15:11]; // extract
  assign n6617_o = n6498_o[20:16]; // extract
  assign n6618_o = n6498_o[22:21]; // extract
  assign n6619_o = n6498_o[23]; // extract
  assign n6620_o = n6498_o[26:24]; // extract
  assign n6621_o = n6498_o[27]; // extract
  assign n6622_o = n6498_o[28]; // extract
  assign n6623_o = n6498_o[29]; // extract
  assign n6624_o = n6498_o[35:30]; // extract
  assign n6625_o = n6498_o[36]; // extract
  assign n6626_o = n6498_o[37]; // extract
  assign n6627_o = n6498_o[38]; // extract
  assign n6628_o = n6498_o[39]; // extract
  assign n6629_o = n6498_o[40]; // extract
  assign n6630_o = n6498_o[43:41]; // extract
  assign n6631_o = n6498_o[55:44]; // extract
  assign n6632_o = n6498_o[62:56]; // extract
  assign n6633_o = n6498_o[63]; // extract
  assign n6634_o = n6498_o[64]; // extract
  assign n6635_o = n6498_o[65]; // extract
  assign n6636_o = n6498_o[66]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:195:24  */
  assign n6637_o = cp_start[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:209:5  */
  neorv32_cpu_cp_muldiv_9159cb8bcee7fcb95582f140960cdae72788d326 neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n6640_o),
    .ctrl_i_rf_rs1(n6641_o),
    .ctrl_i_rf_rs2(n6642_o),
    .ctrl_i_rf_rs3(n6643_o),
    .ctrl_i_rf_rd(n6644_o),
    .ctrl_i_rf_mux(n6645_o),
    .ctrl_i_rf_zero_we(n6646_o),
    .ctrl_i_alu_op(n6647_o),
    .ctrl_i_alu_opa_mux(n6648_o),
    .ctrl_i_alu_opb_mux(n6649_o),
    .ctrl_i_alu_unsigned(n6650_o),
    .ctrl_i_alu_cp_trig(n6651_o),
    .ctrl_i_lsu_req(n6652_o),
    .ctrl_i_lsu_rw(n6653_o),
    .ctrl_i_lsu_mo_we(n6654_o),
    .ctrl_i_lsu_fence(n6655_o),
    .ctrl_i_lsu_priv(n6656_o),
    .ctrl_i_ir_funct3(n6657_o),
    .ctrl_i_ir_funct12(n6658_o),
    .ctrl_i_ir_opcode(n6659_o),
    .ctrl_i_cpu_priv(n6660_o),
    .ctrl_i_cpu_sleep(n6661_o),
    .ctrl_i_cpu_trap(n6662_o),
    .ctrl_i_cpu_debug(n6663_o),
    .start_i(n6664_o),
    .rs1_i(rs1_i),
    .rs2_i(rs2_i),
    .res_o(neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_res_o),
    .valid_o(neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_valid_o));
  assign n6640_o = n6498_o[0]; // extract
  assign n6641_o = n6498_o[5:1]; // extract
  assign n6642_o = n6498_o[10:6]; // extract
  assign n6643_o = n6498_o[15:11]; // extract
  assign n6644_o = n6498_o[20:16]; // extract
  assign n6645_o = n6498_o[22:21]; // extract
  assign n6646_o = n6498_o[23]; // extract
  assign n6647_o = n6498_o[26:24]; // extract
  assign n6648_o = n6498_o[27]; // extract
  assign n6649_o = n6498_o[28]; // extract
  assign n6650_o = n6498_o[29]; // extract
  assign n6651_o = n6498_o[35:30]; // extract
  assign n6652_o = n6498_o[36]; // extract
  assign n6653_o = n6498_o[37]; // extract
  assign n6654_o = n6498_o[38]; // extract
  assign n6655_o = n6498_o[39]; // extract
  assign n6656_o = n6498_o[40]; // extract
  assign n6657_o = n6498_o[43:41]; // extract
  assign n6658_o = n6498_o[55:44]; // extract
  assign n6659_o = n6498_o[62:56]; // extract
  assign n6660_o = n6498_o[63]; // extract
  assign n6661_o = n6498_o[64]; // extract
  assign n6662_o = n6498_o[65]; // extract
  assign n6663_o = n6498_o[66]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_alu.vhd:219:26  */
  assign n6664_o = cp_start[1]; // extract
  assign n6677_o = {n6520_o, n6516_o};
  assign n6678_o = {neorv32_cpu_cp_shifter_inst_res_o, neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_res_o, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  assign n6679_o = {1'b0, 1'b0, 1'b0, 1'b0, neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst_valid_o, neorv32_cpu_cp_shifter_inst_valid_o};
  assign n6686_o = {n6585_o, n6576_o};
endmodule

module neorv32_cpu_regfile_9069ca78e7450a285173431b3e52c5c25299e473
  (input  clk_i,
   input  rstn_i,
   input  ctrl_i_rf_wb_en,
   input  [4:0] ctrl_i_rf_rs1,
   input  [4:0] ctrl_i_rf_rs2,
   input  [4:0] ctrl_i_rf_rs3,
   input  [4:0] ctrl_i_rf_rd,
   input  [1:0] ctrl_i_rf_mux,
   input  ctrl_i_rf_zero_we,
   input  [2:0] ctrl_i_alu_op,
   input  ctrl_i_alu_opa_mux,
   input  ctrl_i_alu_opb_mux,
   input  ctrl_i_alu_unsigned,
   input  [5:0] ctrl_i_alu_cp_trig,
   input  ctrl_i_lsu_req,
   input  ctrl_i_lsu_rw,
   input  ctrl_i_lsu_mo_we,
   input  ctrl_i_lsu_fence,
   input  ctrl_i_lsu_priv,
   input  [2:0] ctrl_i_ir_funct3,
   input  [11:0] ctrl_i_ir_funct12,
   input  [6:0] ctrl_i_ir_opcode,
   input  ctrl_i_cpu_priv,
   input  ctrl_i_cpu_sleep,
   input  ctrl_i_cpu_trap,
   input  ctrl_i_cpu_debug,
   input  [31:0] alu_i,
   input  [31:0] mem_i,
   input  [31:0] csr_i,
   input  [31:0] ret_i,
   output [31:0] rs1_o,
   output [31:0] rs2_o,
   output [31:0] rs3_o,
   output [31:0] rs4_o);
  wire [66:0] n6432_o;
  wire [31:0] rf_wdata;
  wire rf_we;
  wire rd_zero;
  wire [4:0] opa_addr;
  wire [1:0] n6438_o;
  wire n6440_o;
  wire n6442_o;
  wire n6444_o;
  wire n6446_o;
  wire [3:0] n6447_o;
  reg [31:0] n6448_o;
  wire [4:0] n6451_o;
  wire n6453_o;
  wire n6454_o;
  wire n6456_o;
  wire n6457_o;
  wire n6458_o;
  wire n6459_o;
  wire n6460_o;
  wire n6462_o;
  wire [4:0] n6463_o;
  wire [4:0] n6464_o;
  wire n6465_o;
  wire [4:0] n6466_o;
  wire [4:0] n6467_o;
  wire [4:0] n6477_o;
  localparam [31:0] n6485_o = 32'b00000000000000000000000000000000;
  localparam [31:0] n6486_o = 32'b00000000000000000000000000000000;
  reg [31:0] n6494_data; // mem_rd
  reg [31:0] n6496_data; // mem_rd
  assign rs1_o = n6496_data; //(module output)
  assign rs2_o = n6494_data; //(module output)
  assign rs3_o = n6485_o; //(module output)
  assign rs4_o = n6486_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6432_o = {ctrl_i_cpu_debug, ctrl_i_cpu_trap, ctrl_i_cpu_sleep, ctrl_i_cpu_priv, ctrl_i_ir_opcode, ctrl_i_ir_funct12, ctrl_i_ir_funct3, ctrl_i_lsu_priv, ctrl_i_lsu_fence, ctrl_i_lsu_mo_we, ctrl_i_lsu_rw, ctrl_i_lsu_req, ctrl_i_alu_cp_trig, ctrl_i_alu_unsigned, ctrl_i_alu_opb_mux, ctrl_i_alu_opa_mux, ctrl_i_alu_op, ctrl_i_rf_zero_we, ctrl_i_rf_mux, ctrl_i_rf_rd, ctrl_i_rf_rs3, ctrl_i_rf_rs2, ctrl_i_rf_rs1, ctrl_i_rf_wb_en};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:85:10  */
  assign rf_wdata = n6448_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:86:10  */
  assign rf_we = n6460_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:88:10  */
  assign rd_zero = n6454_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:89:10  */
  assign opa_addr = n6463_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:98:17  */
  assign n6438_o = n6432_o[22:21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:99:7  */
  assign n6440_o = n6438_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:100:7  */
  assign n6442_o = n6438_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:101:7  */
  assign n6444_o = n6438_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:102:7  */
  assign n6446_o = n6438_o == 2'b11;
  assign n6447_o = {n6446_o, n6444_o, n6442_o, n6440_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:98:5  */
  always @*
    case (n6447_o)
      4'b1000: n6448_o = ret_i;
      4'b0100: n6448_o = csr_i;
      4'b0010: n6448_o = mem_i;
      4'b0001: n6448_o = alu_i;
      default: n6448_o = alu_i;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:118:34  */
  assign n6451_o = n6432_o[20:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:118:40  */
  assign n6453_o = n6451_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:118:21  */
  assign n6454_o = n6453_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:119:25  */
  assign n6456_o = n6432_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:119:39  */
  assign n6457_o = ~rd_zero;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:119:34  */
  assign n6458_o = n6456_o & n6457_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:119:63  */
  assign n6459_o = n6432_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:119:53  */
  assign n6460_o = n6458_o | n6459_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:120:38  */
  assign n6462_o = n6432_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:120:25  */
  assign n6463_o = n6462_o ? 5'b00000 : n6466_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:121:24  */
  assign n6464_o = n6432_o[20:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:121:43  */
  assign n6465_o = n6432_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:120:56  */
  assign n6466_o = n6465_o ? n6464_o : n6467_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:122:24  */
  assign n6467_o = n6432_o[5:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:131:60  */
  assign n6477_o = n6432_o[10:6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:71:5  */
  reg [31:0] reg_file[31:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n6494_data <= reg_file[n6477_o];
  always @(posedge clk_i)
    if (1'b1)
      n6496_data <= reg_file[opa_addr];
  always @(posedge clk_i)
    if (rf_we)
      reg_file[opa_addr] <= rf_wdata;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:70:5  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:131:26  */
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_regfile.vhd:128:20  */
endmodule

module neorv32_cpu_control_0_64_87d7d7036038d959ad02bd289905a845d3f42491
  (input  clk_i,
   input  clk_aux_i,
   input  rstn_i,
   input  i_pmp_fault_i,
   input  [31:0] bus_rsp_i_data,
   input  bus_rsp_i_ack,
   input  bus_rsp_i_err,
   input  alu_cp_done_i,
   input  [1:0] cmp_i,
   input  [31:0] alu_add_i,
   input  [31:0] rs1_i,
   input  [31:0] xcsr_rdata_i,
   input  db_halt_req_i,
   input  msi_i,
   input  mei_i,
   input  mti_i,
   input  [15:0] firq_i,
   input  lsu_wait_i,
   input  [31:0] mar_i,
   input  ma_load_i,
   input  ma_store_i,
   input  be_load_i,
   input  be_store_i,
   output ctrl_o_rf_wb_en,
   output [4:0] ctrl_o_rf_rs1,
   output [4:0] ctrl_o_rf_rs2,
   output [4:0] ctrl_o_rf_rs3,
   output [4:0] ctrl_o_rf_rd,
   output [1:0] ctrl_o_rf_mux,
   output ctrl_o_rf_zero_we,
   output [2:0] ctrl_o_alu_op,
   output ctrl_o_alu_opa_mux,
   output ctrl_o_alu_opb_mux,
   output ctrl_o_alu_unsigned,
   output [5:0] ctrl_o_alu_cp_trig,
   output ctrl_o_lsu_req,
   output ctrl_o_lsu_rw,
   output ctrl_o_lsu_mo_we,
   output ctrl_o_lsu_fence,
   output ctrl_o_lsu_priv,
   output [2:0] ctrl_o_ir_funct3,
   output [11:0] ctrl_o_ir_funct12,
   output [6:0] ctrl_o_ir_opcode,
   output ctrl_o_cpu_priv,
   output ctrl_o_cpu_sleep,
   output ctrl_o_cpu_trap,
   output ctrl_o_cpu_debug,
   output [31:0] bus_req_o_addr,
   output [31:0] bus_req_o_data,
   output [3:0] bus_req_o_ben,
   output bus_req_o_stb,
   output bus_req_o_rw,
   output bus_req_o_src,
   output bus_req_o_priv,
   output bus_req_o_rvso,
   output bus_req_o_fence,
   output [31:0] imm_o,
   output [31:0] fetch_pc_o,
   output [31:0] curr_pc_o,
   output [31:0] link_pc_o,
   output [31:0] csr_rdata_o,
   output xcsr_we_o,
   output [11:0] xcsr_addr_o,
   output [31:0] xcsr_wdata_o);
  wire n2328_o;
  wire [4:0] n2329_o;
  wire [4:0] n2330_o;
  wire [4:0] n2331_o;
  wire [4:0] n2332_o;
  wire [1:0] n2333_o;
  wire n2334_o;
  wire [2:0] n2335_o;
  wire n2336_o;
  wire n2337_o;
  wire n2338_o;
  wire [5:0] n2339_o;
  wire n2340_o;
  wire n2341_o;
  wire n2342_o;
  wire n2343_o;
  wire n2344_o;
  wire [2:0] n2345_o;
  wire [11:0] n2346_o;
  wire [6:0] n2347_o;
  wire n2348_o;
  wire n2349_o;
  wire n2350_o;
  wire n2351_o;
  wire [31:0] n2353_o;
  wire [31:0] n2354_o;
  wire [3:0] n2355_o;
  wire n2356_o;
  wire n2357_o;
  wire n2358_o;
  wire n2359_o;
  wire n2360_o;
  wire n2361_o;
  wire [33:0] n2362_o;
  wire [37:0] fetch_engine;
  wire [75:0] ipb;
  wire [87:0] issue_engine;
  wire [16:0] decode_aux;
  wire [203:0] execute_engine;
  wire [20:0] monitor;
  wire sleep_mode;
  wire [103:0] trap_ctrl;
  wire [66:0] ctrl;
  wire [66:0] ctrl_nxt;
  wire [507:0] csr;
  wire [341:0] cnt;
  wire [95:0] cnt_lo_rd;
  wire [95:0] cnt_hi_rd;
  wire [11:0] cnt_event;
  wire [4:0] debug_ctrl;
  wire illegal_cmd;
  wire csr_reg_valid;
  wire csr_rw_valid;
  wire csr_priv_valid;
  wire hw_trigger_fired;
  wire [31:0] csr_rdata;
  wire [31:0] xcsr_rdata;
  wire n2372_o;
  wire [1:0] n2378_o;
  wire n2380_o;
  wire n2382_o;
  wire n2383_o;
  wire n2384_o;
  wire n2385_o;
  wire [1:0] n2386_o;
  wire [1:0] n2387_o;
  wire n2389_o;
  wire n2391_o;
  wire n2392_o;
  wire n2393_o;
  wire [1:0] n2395_o;
  wire [1:0] n2396_o;
  wire [1:0] n2397_o;
  wire n2399_o;
  wire n2400_o;
  wire [31:0] n2401_o;
  wire [31:0] n2403_o;
  wire [29:0] n2405_o;
  wire n2406_o;
  wire n2407_o;
  wire n2408_o;
  wire n2409_o;
  wire [1:0] n2412_o;
  wire [31:0] n2413_o;
  wire [1:0] n2414_o;
  wire [1:0] n2415_o;
  wire [31:0] n2416_o;
  wire [31:0] n2417_o;
  wire n2419_o;
  wire [30:0] n2420_o;
  wire [31:0] n2422_o;
  wire n2423_o;
  wire [1:0] n2425_o;
  reg [1:0] n2426_o;
  wire [31:0] n2427_o;
  reg [31:0] n2428_o;
  wire n2429_o;
  reg n2430_o;
  wire [34:0] n2431_o;
  wire [34:0] n2436_o;
  wire [29:0] n2440_o;
  wire [31:0] n2442_o;
  wire [29:0] n2443_o;
  wire [31:0] n2445_o;
  wire [1:0] n2447_o;
  wire n2449_o;
  wire [1:0] n2450_o;
  wire n2452_o;
  wire n2453_o;
  wire n2454_o;
  wire n2456_o;
  wire n2457_o;
  wire n2458_o;
  wire n2459_o;
  wire n2460_o;
  wire [15:0] n2461_o;
  wire [16:0] n2462_o;
  wire n2463_o;
  wire n2464_o;
  wire [15:0] n2465_o;
  wire [16:0] n2466_o;
  wire [1:0] n2468_o;
  wire n2470_o;
  wire n2471_o;
  wire n2472_o;
  wire n2473_o;
  wire n2474_o;
  wire n2476_o;
  wire n2477_o;
  wire n2478_o;
  wire [1:0] n2481_o;
  wire n2483_o;
  wire n2484_o;
  wire n2485_o;
  wire n2486_o;
  wire n2488_o;
  wire n2494_o;
  wire prefetch_buffer_n1_prefetch_buffer_inst_half_o;
  wire prefetch_buffer_n1_prefetch_buffer_inst_free_o;
  wire [16:0] prefetch_buffer_n1_prefetch_buffer_inst_rdata_o;
  wire prefetch_buffer_n1_prefetch_buffer_inst_avail_o;
  wire n2495_o;
  wire [16:0] n2496_o;
  wire n2497_o;
  wire n2499_o;
  wire prefetch_buffer_n2_prefetch_buffer_inst_half_o;
  wire prefetch_buffer_n2_prefetch_buffer_inst_free_o;
  wire [16:0] prefetch_buffer_n2_prefetch_buffer_inst_rdata_o;
  wire prefetch_buffer_n2_prefetch_buffer_inst_avail_o;
  wire n2502_o;
  wire [16:0] n2503_o;
  wire n2504_o;
  wire n2506_o;
  wire [31:0] neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_instr32_o;
  wire [15:0] n2509_o;
  wire [15:0] n2511_o;
  wire n2512_o;
  wire n2513_o;
  wire [15:0] n2514_o;
  wire [15:0] n2515_o;
  wire n2517_o;
  wire n2520_o;
  wire n2521_o;
  wire n2522_o;
  wire n2523_o;
  wire n2524_o;
  wire n2525_o;
  wire n2526_o;
  wire n2527_o;
  wire n2528_o;
  wire n2529_o;
  wire n2530_o;
  wire n2531_o;
  localparam [1:0] n2539_o = 2'b00;
  wire n2540_o;
  wire n2541_o;
  wire [1:0] n2542_o;
  wire n2544_o;
  wire n2545_o;
  wire n2546_o;
  wire n2547_o;
  wire [1:0] n2549_o;
  wire [31:0] n2550_o;
  wire [33:0] n2551_o;
  wire n2552_o;
  wire n2553_o;
  wire n2554_o;
  wire n2555_o;
  wire n2556_o;
  wire n2557_o;
  wire [1:0] n2558_o;
  wire n2559_o;
  wire [1:0] n2561_o;
  wire [15:0] n2562_o;
  wire [17:0] n2563_o;
  wire [15:0] n2564_o;
  wire [33:0] n2565_o;
  wire [35:0] n2566_o;
  wire [34:0] n2567_o;
  wire n2568_o;
  wire [34:0] n2569_o;
  wire [34:0] n2570_o;
  wire n2571_o;
  wire n2572_o;
  wire n2573_o;
  wire [1:0] n2574_o;
  wire n2576_o;
  wire n2577_o;
  wire n2578_o;
  wire n2579_o;
  wire [1:0] n2581_o;
  wire [31:0] n2582_o;
  wire [33:0] n2583_o;
  wire n2584_o;
  wire n2585_o;
  wire n2586_o;
  wire n2587_o;
  wire n2588_o;
  wire n2589_o;
  wire [1:0] n2590_o;
  wire n2591_o;
  wire [1:0] n2593_o;
  wire [15:0] n2594_o;
  wire [17:0] n2595_o;
  wire [15:0] n2596_o;
  wire [33:0] n2597_o;
  wire [35:0] n2598_o;
  wire n2599_o;
  wire [33:0] n2600_o;
  wire [33:0] n2601_o;
  wire n2602_o;
  wire n2603_o;
  wire n2604_o;
  wire n2605_o;
  wire n2606_o;
  wire [35:0] n2607_o;
  wire [35:0] n2608_o;
  wire n2609_o;
  wire n2610_o;
  wire [35:0] n2611_o;
  wire n2613_o;
  wire n2614_o;
  wire n2615_o;
  wire n2616_o;
  wire n2617_o;
  wire n2618_o;
  wire n2620_o;
  wire n2622_o;
  wire n2623_o;
  wire n2624_o;
  wire n2625_o;
  wire n2626_o;
  wire n2627_o;
  wire n2628_o;
  wire n2629_o;
  wire n2630_o;
  wire n2631_o;
  wire n2632_o;
  wire n2633_o;
  wire n2634_o;
  wire n2635_o;
  wire n2636_o;
  wire n2637_o;
  wire n2638_o;
  wire n2639_o;
  wire n2640_o;
  wire n2641_o;
  wire n2642_o;
  wire [3:0] n2643_o;
  wire [3:0] n2644_o;
  wire [3:0] n2645_o;
  wire [3:0] n2646_o;
  wire [3:0] n2647_o;
  wire [15:0] n2648_o;
  wire [4:0] n2649_o;
  wire [20:0] n2650_o;
  wire n2652_o;
  wire [6:0] n2653_o;
  wire n2654_o;
  wire n2655_o;
  wire n2656_o;
  wire n2657_o;
  wire n2658_o;
  wire n2659_o;
  wire n2660_o;
  wire n2661_o;
  wire n2662_o;
  wire n2663_o;
  wire n2664_o;
  wire n2665_o;
  wire n2666_o;
  wire n2667_o;
  wire n2668_o;
  wire n2669_o;
  wire n2670_o;
  wire n2671_o;
  wire n2672_o;
  wire n2673_o;
  wire n2674_o;
  wire [3:0] n2675_o;
  wire [3:0] n2676_o;
  wire [3:0] n2677_o;
  wire [3:0] n2678_o;
  wire [3:0] n2679_o;
  wire [15:0] n2680_o;
  wire [4:0] n2681_o;
  wire [20:0] n2682_o;
  wire [5:0] n2683_o;
  wire [4:0] n2684_o;
  wire n2686_o;
  wire n2687_o;
  wire n2688_o;
  wire n2689_o;
  wire n2690_o;
  wire n2691_o;
  wire n2692_o;
  wire n2693_o;
  wire n2694_o;
  wire n2695_o;
  wire n2696_o;
  wire n2697_o;
  wire n2698_o;
  wire n2699_o;
  wire n2700_o;
  wire n2701_o;
  wire n2702_o;
  wire n2703_o;
  wire n2704_o;
  wire n2705_o;
  wire n2706_o;
  wire [3:0] n2707_o;
  wire [3:0] n2708_o;
  wire [3:0] n2709_o;
  wire [3:0] n2710_o;
  wire [3:0] n2711_o;
  wire [15:0] n2712_o;
  wire [19:0] n2713_o;
  wire n2714_o;
  wire [5:0] n2715_o;
  wire [3:0] n2716_o;
  wire n2719_o;
  wire [19:0] n2720_o;
  localparam [11:0] n2721_o = 12'b000000000000;
  wire n2723_o;
  wire n2725_o;
  wire n2726_o;
  wire n2727_o;
  wire n2728_o;
  wire n2729_o;
  wire n2730_o;
  wire n2731_o;
  wire n2732_o;
  wire n2733_o;
  wire n2734_o;
  wire n2735_o;
  wire n2736_o;
  wire n2737_o;
  wire n2738_o;
  wire [3:0] n2739_o;
  wire [3:0] n2740_o;
  wire [3:0] n2741_o;
  wire [11:0] n2742_o;
  wire [7:0] n2743_o;
  wire n2744_o;
  wire [9:0] n2745_o;
  wire n2748_o;
  wire n2750_o;
  wire [4:0] n2751_o;
  wire n2752_o;
  wire n2753_o;
  reg n2754_o;
  wire [3:0] n2755_o;
  wire [3:0] n2756_o;
  wire [3:0] n2757_o;
  wire [3:0] n2758_o;
  reg [3:0] n2759_o;
  wire [5:0] n2760_o;
  wire [5:0] n2761_o;
  wire [5:0] n2762_o;
  reg [5:0] n2763_o;
  wire n2764_o;
  wire n2765_o;
  wire n2766_o;
  reg n2767_o;
  wire [7:0] n2768_o;
  wire [7:0] n2769_o;
  wire [7:0] n2770_o;
  wire [7:0] n2771_o;
  reg [7:0] n2772_o;
  wire [11:0] n2773_o;
  wire [11:0] n2774_o;
  wire [11:0] n2775_o;
  wire [11:0] n2776_o;
  reg [11:0] n2777_o;
  wire [31:0] n2781_o;
  wire n2787_o;
  wire n2788_o;
  wire n2789_o;
  wire n2790_o;
  wire n2791_o;
  wire n2792_o;
  wire n2793_o;
  wire n2794_o;
  wire n2795_o;
  wire n2796_o;
  wire n2797_o;
  wire n2799_o;
  wire n2802_o;
  wire [3:0] n2810_o;
  wire [31:0] n2811_o;
  wire n2812_o;
  wire n2813_o;
  wire [30:0] n2814_o;
  wire [31:0] n2816_o;
  wire [3:0] n2819_o;
  wire n2821_o;
  wire [30:0] n2822_o;
  wire [31:0] n2824_o;
  wire [3:0] n2827_o;
  wire [1:0] n2830_o;
  wire n2832_o;
  wire n2833_o;
  wire n2834_o;
  wire [24:0] n2835_o;
  wire [4:0] n2836_o;
  wire [29:0] n2837_o;
  wire [31:0] n2839_o;
  wire [29:0] n2840_o;
  wire [31:0] n2842_o;
  wire [31:0] n2843_o;
  wire n2845_o;
  wire [30:0] n2847_o;
  wire [31:0] n2849_o;
  wire n2851_o;
  wire n2852_o;
  wire n2853_o;
  wire n2854_o;
  wire n2855_o;
  wire [30:0] n2856_o;
  wire [31:0] n2858_o;
  wire [31:0] n2859_o;
  wire [31:0] n2860_o;
  wire n2862_o;
  wire [31:0] n2863_o;
  wire [31:0] n2864_o;
  wire [31:0] n2865_o;
  wire n2867_o;
  wire [3:0] n2868_o;
  wire [31:0] n2869_o;
  reg [31:0] n2870_o;
  wire n2905_o;
  wire n2909_o;
  wire n2910_o;
  wire n2912_o;
  wire [3:0] n2913_o;
  wire [30:0] n2915_o;
  wire [31:0] n2917_o;
  wire [30:0] n2918_o;
  wire [31:0] n2920_o;
  wire [6:0] n2930_o;
  wire n2932_o;
  wire n2933_o;
  wire n2934_o;
  wire n2936_o;
  wire n2938_o;
  wire n2939_o;
  wire n2941_o;
  wire n2943_o;
  wire [1:0] n2944_o;
  wire [1:0] n2945_o;
  wire [1:0] n2946_o;
  wire [4:0] n2949_o;
  wire n2951_o;
  wire n2952_o;
  wire [4:0] n2955_o;
  wire n2957_o;
  wire n2958_o;
  wire [4:0] n2960_o;
  wire [6:0] n2962_o;
  wire [3:0] n2964_o;
  wire [31:0] n2965_o;
  wire n2966_o;
  wire n2978_o;
  wire n2979_o;
  wire n2980_o;
  wire n2981_o;
  localparam [66:0] n2982_o = 67'b0000000000000000000000000000000000000000000000000000000000000000000;
  wire [6:0] n2985_o;
  wire n2988_o;
  wire n2990_o;
  wire n2991_o;
  wire n2993_o;
  wire n2994_o;
  reg n2996_o;
  wire [6:0] n2999_o;
  wire n3002_o;
  wire n3004_o;
  wire n3005_o;
  wire n3007_o;
  wire n3008_o;
  wire n3010_o;
  wire n3011_o;
  wire n3013_o;
  wire n3014_o;
  wire n3016_o;
  wire n3017_o;
  wire n3019_o;
  wire n3020_o;
  wire n3022_o;
  wire n3023_o;
  wire n3025_o;
  wire n3026_o;
  reg n3028_o;
  wire n3029_o;
  wire [3:0] n3032_o;
  wire n3033_o;
  wire n3034_o;
  wire n3035_o;
  wire n3037_o;
  wire n3038_o;
  wire n3039_o;
  wire n3041_o;
  wire n3042_o;
  wire [31:0] n3043_o;
  wire n3046_o;
  wire [3:0] n3047_o;
  wire [31:0] n3048_o;
  wire n3049_o;
  wire n3050_o;
  wire n3051_o;
  wire n3052_o;
  wire [3:0] n3053_o;
  wire [31:0] n3054_o;
  wire n3055_o;
  wire n3056_o;
  wire n3057_o;
  wire n3059_o;
  wire n3060_o;
  wire [3:0] n3063_o;
  wire n3064_o;
  wire n3066_o;
  wire n3070_o;
  wire n3074_o;
  wire [6:0] n3075_o;
  wire [2:0] n3076_o;
  wire n3077_o;
  wire n3078_o;
  wire n3079_o;
  wire [2:0] n3082_o;
  wire n3084_o;
  wire n3087_o;
  wire n3089_o;
  wire n3090_o;
  wire n3093_o;
  wire n3096_o;
  wire [3:0] n3098_o;
  reg [2:0] n3099_o;
  wire n3100_o;
  wire n3102_o;
  wire n3103_o;
  wire n3104_o;
  wire n3105_o;
  wire n3106_o;
  wire n3108_o;
  wire [2:0] n3111_o;
  wire n3113_o;
  wire [2:0] n3114_o;
  wire n3116_o;
  wire n3117_o;
  wire [3:0] n3122_o;
  wire n3123_o;
  wire n3124_o;
  wire n3125_o;
  wire n3126_o;
  wire [3:0] n3127_o;
  wire n3128_o;
  wire n3129_o;
  wire n3130_o;
  wire n3131_o;
  wire n3132_o;
  wire n3133_o;
  wire n3135_o;
  wire n3137_o;
  wire n3138_o;
  wire n3139_o;
  wire [2:0] n3141_o;
  wire n3145_o;
  wire n3147_o;
  wire n3148_o;
  wire n3151_o;
  wire n3153_o;
  wire n3154_o;
  wire n3156_o;
  wire n3157_o;
  wire n3160_o;
  wire n3162_o;
  wire n3163_o;
  wire n3165_o;
  wire n3166_o;
  wire n3169_o;
  wire n3173_o;
  wire n3177_o;
  wire n3179_o;
  wire n3180_o;
  wire n3182_o;
  wire n3183_o;
  wire n3185_o;
  wire n3186_o;
  wire [6:0] n3189_o;
  reg [3:0] n3190_o;
  wire n3191_o;
  reg n3192_o;
  wire [2:0] n3193_o;
  reg [2:0] n3194_o;
  wire n3195_o;
  reg n3196_o;
  wire n3197_o;
  reg n3198_o;
  wire n3199_o;
  reg n3200_o;
  wire n3201_o;
  reg n3202_o;
  reg n3203_o;
  wire n3205_o;
  wire n3207_o;
  wire n3208_o;
  wire [3:0] n3211_o;
  wire n3212_o;
  wire n3213_o;
  wire n3215_o;
  wire n3216_o;
  wire [3:0] n3220_o;
  wire n3221_o;
  wire n3222_o;
  wire n3224_o;
  wire n3226_o;
  wire n3227_o;
  wire n3228_o;
  wire n3229_o;
  wire n3230_o;
  wire n3234_o;
  wire [3:0] n3235_o;
  wire n3237_o;
  wire n3242_o;
  wire n3243_o;
  wire [3:0] n3247_o;
  wire n3248_o;
  wire n3249_o;
  wire n3251_o;
  wire n3253_o;
  wire n3254_o;
  wire n3255_o;
  wire n3256_o;
  wire n3257_o;
  wire n3258_o;
  wire n3259_o;
  wire n3260_o;
  wire n3261_o;
  wire n3262_o;
  wire n3263_o;
  wire n3265_o;
  wire n3267_o;
  wire n3268_o;
  wire [3:0] n3270_o;
  wire n3272_o;
  wire n3274_o;
  wire n3275_o;
  wire [3:0] n3277_o;
  wire n3279_o;
  wire [2:0] n3281_o;
  wire n3283_o;
  wire n3284_o;
  wire n3285_o;
  wire n3286_o;
  wire [11:0] n3287_o;
  wire n3290_o;
  wire n3293_o;
  wire n3296_o;
  wire n3298_o;
  wire n3299_o;
  wire [2:0] n3301_o;
  reg [3:0] n3302_o;
  reg n3303_o;
  reg n3304_o;
  wire [2:0] n3305_o;
  wire n3307_o;
  wire [2:0] n3308_o;
  wire n3310_o;
  wire n3311_o;
  wire n3312_o;
  wire n3313_o;
  wire n3314_o;
  wire n3316_o;
  wire [3:0] n3318_o;
  wire [1:0] n3319_o;
  wire [1:0] n3320_o;
  wire [1:0] n3321_o;
  wire n3322_o;
  wire n3323_o;
  wire n3324_o;
  wire [11:0] n3325_o;
  reg n3326_o;
  reg n3327_o;
  reg [3:0] n3328_o;
  reg [31:0] n3329_o;
  reg n3330_o;
  reg n3331_o;
  reg n3332_o;
  reg n3333_o;
  reg n3334_o;
  wire [1:0] n3335_o;
  reg [1:0] n3336_o;
  wire n3337_o;
  reg n3338_o;
  wire [1:0] n3339_o;
  reg [1:0] n3340_o;
  wire n3341_o;
  reg n3342_o;
  wire [2:0] n3343_o;
  reg [2:0] n3344_o;
  wire n3345_o;
  reg n3346_o;
  wire n3347_o;
  reg n3348_o;
  wire n3349_o;
  reg n3350_o;
  wire n3351_o;
  reg n3352_o;
  wire n3353_o;
  reg n3354_o;
  wire n3355_o;
  reg n3356_o;
  wire [19:0] n3359_o;
  wire n3364_o;
  wire n3366_o;
  wire [26:0] n3367_o;
  wire n3368_o;
  reg n3369_o;
  reg n3370_o;
  wire n3373_o;
  wire [3:0] n3375_o;
  wire n3377_o;
  wire [1:0] n3378_o;
  wire n3380_o;
  wire n3381_o;
  wire n3382_o;
  wire n3383_o;
  wire n3384_o;
  wire n3387_o;
  wire n3392_o;
  wire n3393_o;
  wire n3394_o;
  wire n3395_o;
  wire n3396_o;
  wire n3397_o;
  wire n3398_o;
  wire n3399_o;
  wire n3400_o;
  wire n3401_o;
  wire n3402_o;
  wire n3403_o;
  wire n3404_o;
  wire n3405_o;
  wire n3406_o;
  wire n3407_o;
  wire n3408_o;
  wire n3409_o;
  wire n3410_o;
  wire n3411_o;
  wire n3412_o;
  wire n3413_o;
  wire [4:0] n3414_o;
  wire [4:0] n3415_o;
  wire [4:0] n3416_o;
  wire [4:0] n3417_o;
  wire [1:0] n3418_o;
  wire n3419_o;
  wire [2:0] n3420_o;
  wire n3421_o;
  wire n3422_o;
  wire n3423_o;
  wire [5:0] n3424_o;
  wire n3425_o;
  wire n3426_o;
  wire [3:0] n3428_o;
  wire n3430_o;
  wire n3431_o;
  wire n3433_o;
  wire n3434_o;
  wire n3435_o;
  wire n3436_o;
  wire n3437_o;
  wire [2:0] n3438_o;
  wire [11:0] n3439_o;
  wire [6:0] n3440_o;
  wire n3441_o;
  wire n3442_o;
  wire n3443_o;
  wire n3445_o;
  wire [9:0] n3448_o;
  wire [9:0] n3450_o;
  wire [9:0] n3455_o;
  wire [3:0] n3456_o;
  wire n3458_o;
  wire [9:0] n3459_o;
  wire n3461_o;
  wire [11:0] n3463_o;
  wire n3466_o;
  wire n3468_o;
  wire n3469_o;
  wire n3471_o;
  wire n3472_o;
  wire n3474_o;
  wire n3475_o;
  wire n3478_o;
  wire n3480_o;
  wire n3481_o;
  wire n3483_o;
  wire n3484_o;
  wire n3486_o;
  wire n3488_o;
  wire n3489_o;
  wire n3491_o;
  wire n3492_o;
  wire n3494_o;
  wire n3495_o;
  wire n3497_o;
  wire n3498_o;
  wire n3500_o;
  wire n3501_o;
  wire n3503_o;
  wire n3504_o;
  wire n3506_o;
  wire n3507_o;
  wire n3509_o;
  wire n3510_o;
  wire n3512_o;
  wire n3513_o;
  wire n3515_o;
  wire n3516_o;
  wire n3518_o;
  wire n3519_o;
  wire n3521_o;
  wire n3522_o;
  wire n3524_o;
  wire n3525_o;
  wire n3527_o;
  wire n3528_o;
  wire n3530_o;
  wire n3531_o;
  wire n3533_o;
  wire n3534_o;
  wire n3536_o;
  wire n3537_o;
  wire n3540_o;
  wire n3542_o;
  wire n3543_o;
  wire n3545_o;
  wire n3546_o;
  wire n3549_o;
  wire n3551_o;
  wire n3552_o;
  wire n3554_o;
  wire n3555_o;
  wire n3557_o;
  wire n3558_o;
  wire n3560_o;
  wire n3561_o;
  wire n3563_o;
  wire n3564_o;
  wire n3566_o;
  wire n3567_o;
  wire n3569_o;
  wire n3570_o;
  wire n3572_o;
  wire n3573_o;
  wire n3575_o;
  wire n3576_o;
  wire n3578_o;
  wire n3579_o;
  wire n3581_o;
  wire n3582_o;
  wire n3584_o;
  wire n3585_o;
  wire n3587_o;
  wire n3588_o;
  wire n3590_o;
  wire n3591_o;
  wire n3593_o;
  wire n3594_o;
  wire n3596_o;
  wire n3597_o;
  wire n3599_o;
  wire n3600_o;
  wire n3602_o;
  wire n3603_o;
  wire n3605_o;
  wire n3606_o;
  wire n3609_o;
  wire n3611_o;
  wire n3612_o;
  wire n3614_o;
  wire n3615_o;
  wire n3617_o;
  wire n3618_o;
  wire n3620_o;
  wire n3621_o;
  wire n3623_o;
  wire n3624_o;
  wire n3626_o;
  wire n3627_o;
  wire n3629_o;
  wire n3630_o;
  wire n3632_o;
  wire n3633_o;
  wire n3635_o;
  wire n3636_o;
  wire n3638_o;
  wire n3639_o;
  wire n3641_o;
  wire n3642_o;
  wire n3644_o;
  wire n3645_o;
  wire n3647_o;
  wire n3648_o;
  wire n3650_o;
  wire n3651_o;
  wire n3653_o;
  wire n3654_o;
  wire n3656_o;
  wire n3657_o;
  wire n3659_o;
  wire n3660_o;
  wire n3662_o;
  wire n3663_o;
  wire n3665_o;
  wire n3666_o;
  wire n3668_o;
  wire n3669_o;
  wire n3671_o;
  wire n3672_o;
  wire n3674_o;
  wire n3675_o;
  wire n3677_o;
  wire n3678_o;
  wire n3680_o;
  wire n3681_o;
  wire n3683_o;
  wire n3684_o;
  wire n3686_o;
  wire n3687_o;
  wire n3689_o;
  wire n3690_o;
  wire n3692_o;
  wire n3693_o;
  wire n3695_o;
  wire n3696_o;
  wire n3698_o;
  wire n3699_o;
  wire n3701_o;
  wire n3702_o;
  wire n3704_o;
  wire n3705_o;
  wire n3707_o;
  wire n3708_o;
  wire n3710_o;
  wire n3711_o;
  wire n3713_o;
  wire n3714_o;
  wire n3716_o;
  wire n3717_o;
  wire n3719_o;
  wire n3720_o;
  wire n3722_o;
  wire n3723_o;
  wire n3725_o;
  wire n3726_o;
  wire n3728_o;
  wire n3729_o;
  wire n3731_o;
  wire n3732_o;
  wire n3734_o;
  wire n3735_o;
  wire n3737_o;
  wire n3738_o;
  wire n3740_o;
  wire n3741_o;
  wire n3743_o;
  wire n3744_o;
  wire n3746_o;
  wire n3747_o;
  wire n3749_o;
  wire n3750_o;
  wire n3752_o;
  wire n3753_o;
  wire n3755_o;
  wire n3756_o;
  wire n3758_o;
  wire n3759_o;
  wire n3761_o;
  wire n3762_o;
  wire n3764_o;
  wire n3765_o;
  wire n3767_o;
  wire n3768_o;
  wire n3770_o;
  wire n3771_o;
  wire n3773_o;
  wire n3774_o;
  wire n3776_o;
  wire n3777_o;
  wire n3779_o;
  wire n3780_o;
  wire n3782_o;
  wire n3783_o;
  wire n3785_o;
  wire n3786_o;
  wire n3788_o;
  wire n3789_o;
  wire n3791_o;
  wire n3792_o;
  wire n3794_o;
  wire n3795_o;
  wire n3797_o;
  wire n3798_o;
  wire n3800_o;
  wire n3801_o;
  wire n3804_o;
  wire n3806_o;
  wire n3807_o;
  wire n3809_o;
  wire n3810_o;
  wire n3812_o;
  wire n3813_o;
  wire n3815_o;
  wire n3816_o;
  wire n3818_o;
  wire n3819_o;
  wire n3821_o;
  wire n3822_o;
  wire n3824_o;
  wire n3825_o;
  wire n3828_o;
  wire n3830_o;
  wire n3831_o;
  wire n3833_o;
  wire n3834_o;
  wire n3837_o;
  wire n3839_o;
  wire n3840_o;
  wire n3842_o;
  wire n3843_o;
  wire n3845_o;
  wire n3846_o;
  wire [8:0] n3847_o;
  reg n3858_o;
  wire [1:0] n3861_o;
  wire n3863_o;
  wire [2:0] n3864_o;
  wire n3866_o;
  wire [2:0] n3867_o;
  wire n3869_o;
  wire n3870_o;
  wire n3871_o;
  wire n3872_o;
  wire n3873_o;
  wire n3874_o;
  wire n3877_o;
  wire [3:0] n3891_o;
  wire n3893_o;
  wire n3895_o;
  wire n3897_o;
  wire n3898_o;
  wire n3899_o;
  wire n3900_o;
  wire n3901_o;
  wire n3902_o;
  wire n3903_o;
  wire [1:0] n3904_o;
  wire n3906_o;
  wire n3907_o;
  wire n3908_o;
  wire n3909_o;
  wire n3912_o;
  wire n3914_o;
  wire [6:0] n3917_o;
  wire n3919_o;
  wire n3921_o;
  wire n3922_o;
  wire n3924_o;
  wire n3925_o;
  wire [2:0] n3926_o;
  wire n3928_o;
  reg n3931_o;
  wire n3933_o;
  wire [2:0] n3934_o;
  wire n3936_o;
  wire n3938_o;
  wire n3939_o;
  wire n3941_o;
  wire n3942_o;
  wire n3944_o;
  wire n3945_o;
  wire n3947_o;
  wire n3948_o;
  wire n3950_o;
  wire n3951_o;
  reg n3954_o;
  wire n3956_o;
  wire [2:0] n3957_o;
  wire n3959_o;
  wire n3961_o;
  wire n3962_o;
  wire n3964_o;
  wire n3965_o;
  wire n3967_o;
  wire n3968_o;
  wire n3970_o;
  wire n3971_o;
  reg n3974_o;
  wire n3976_o;
  wire [2:0] n3977_o;
  wire n3979_o;
  wire n3981_o;
  wire n3982_o;
  wire n3984_o;
  wire n3985_o;
  reg n3988_o;
  wire n3990_o;
  wire n3992_o;
  wire [2:0] n3993_o;
  wire n3995_o;
  wire [2:0] n3996_o;
  wire n3998_o;
  wire n3999_o;
  wire [4:0] n4000_o;
  wire n4002_o;
  wire n4003_o;
  wire n4004_o;
  wire n4005_o;
  wire n4006_o;
  wire [2:0] n4007_o;
  wire n4009_o;
  wire [2:0] n4010_o;
  wire n4012_o;
  wire n4013_o;
  wire [2:0] n4014_o;
  wire n4016_o;
  wire n4017_o;
  wire [2:0] n4018_o;
  wire n4020_o;
  wire n4021_o;
  wire [2:0] n4022_o;
  wire n4024_o;
  wire n4025_o;
  wire [2:0] n4026_o;
  wire n4028_o;
  wire n4029_o;
  wire [6:0] n4030_o;
  wire n4032_o;
  wire n4033_o;
  wire n4034_o;
  wire n4035_o;
  wire n4037_o;
  wire n4038_o;
  wire n4039_o;
  wire n4041_o;
  wire n4042_o;
  wire n4044_o;
  wire n4046_o;
  wire n4049_o;
  wire n4051_o;
  wire [2:0] n4052_o;
  wire n4054_o;
  wire [2:0] n4055_o;
  wire n4057_o;
  wire n4058_o;
  wire [2:0] n4059_o;
  wire n4061_o;
  wire n4062_o;
  wire [2:0] n4063_o;
  wire n4065_o;
  wire n4066_o;
  wire [2:0] n4067_o;
  wire n4069_o;
  wire n4070_o;
  wire [2:0] n4071_o;
  wire n4073_o;
  wire n4074_o;
  wire [2:0] n4075_o;
  wire n4077_o;
  wire [6:0] n4078_o;
  wire n4080_o;
  wire n4081_o;
  wire n4082_o;
  wire [2:0] n4083_o;
  wire n4085_o;
  wire [4:0] n4086_o;
  wire n4088_o;
  wire n4089_o;
  wire n4090_o;
  wire n4091_o;
  wire n4092_o;
  wire n4093_o;
  wire n4095_o;
  wire n4098_o;
  wire n4100_o;
  wire [2:0] n4101_o;
  wire n4103_o;
  wire n4105_o;
  wire n4106_o;
  reg n4109_o;
  wire n4111_o;
  wire [2:0] n4112_o;
  wire n4114_o;
  wire n4115_o;
  wire n4116_o;
  wire n4117_o;
  wire [11:0] n4118_o;
  wire n4120_o;
  wire n4122_o;
  wire n4123_o;
  wire n4124_o;
  wire n4125_o;
  wire n4126_o;
  wire n4127_o;
  wire n4129_o;
  wire n4130_o;
  wire n4131_o;
  wire n4133_o;
  wire n4134_o;
  wire n4135_o;
  wire n4136_o;
  wire n4137_o;
  wire n4139_o;
  wire [3:0] n4140_o;
  reg n4143_o;
  wire n4145_o;
  wire n4146_o;
  wire n4147_o;
  wire n4148_o;
  wire n4149_o;
  wire n4150_o;
  wire [2:0] n4151_o;
  wire n4153_o;
  wire n4154_o;
  wire n4157_o;
  wire n4158_o;
  wire n4160_o;
  wire n4162_o;
  wire n4163_o;
  wire n4165_o;
  wire n4167_o;
  wire n4170_o;
  wire n4172_o;
  wire n4173_o;
  wire n4175_o;
  wire n4176_o;
  wire n4178_o;
  wire n4179_o;
  wire [11:0] n4180_o;
  reg n4185_o;
  wire [3:0] n4189_o;
  wire n4191_o;
  wire [3:0] n4192_o;
  wire n4194_o;
  wire n4195_o;
  wire n4196_o;
  wire n4197_o;
  wire [1:0] n4198_o;
  wire n4200_o;
  wire n4201_o;
  wire n4202_o;
  wire n4203_o;
  wire n4206_o;
  wire n4209_o;
  wire n4210_o;
  wire n4211_o;
  wire n4212_o;
  wire n4213_o;
  wire n4214_o;
  wire n4215_o;
  wire n4216_o;
  wire n4217_o;
  wire n4218_o;
  wire n4219_o;
  wire n4220_o;
  wire n4221_o;
  wire n4222_o;
  wire n4223_o;
  wire n4224_o;
  wire n4225_o;
  wire n4226_o;
  wire n4227_o;
  wire n4228_o;
  wire n4229_o;
  wire n4230_o;
  wire n4231_o;
  wire n4232_o;
  wire n4233_o;
  wire n4234_o;
  wire n4235_o;
  wire n4236_o;
  wire n4237_o;
  wire n4238_o;
  wire n4239_o;
  wire n4240_o;
  wire n4241_o;
  wire n4242_o;
  wire n4243_o;
  wire n4244_o;
  wire n4245_o;
  wire n4246_o;
  wire n4247_o;
  wire n4248_o;
  wire n4249_o;
  wire n4250_o;
  wire n4251_o;
  wire n4252_o;
  wire n4253_o;
  wire n4254_o;
  wire n4255_o;
  wire n4256_o;
  wire n4257_o;
  wire n4258_o;
  wire n4259_o;
  wire n4260_o;
  wire n4261_o;
  wire n4262_o;
  wire n4263_o;
  wire [10:0] n4266_o;
  wire n4272_o;
  wire n4276_o;
  wire n4278_o;
  wire n4279_o;
  wire n4280_o;
  wire n4281_o;
  wire n4283_o;
  wire n4284_o;
  wire n4285_o;
  wire n4286_o;
  wire n4288_o;
  wire n4289_o;
  wire n4290_o;
  wire n4291_o;
  wire n4293_o;
  wire n4294_o;
  wire n4295_o;
  wire n4296_o;
  wire n4298_o;
  wire n4299_o;
  wire n4300_o;
  wire n4301_o;
  wire n4303_o;
  wire n4304_o;
  wire n4305_o;
  wire n4306_o;
  wire n4308_o;
  wire n4309_o;
  wire n4310_o;
  wire n4311_o;
  wire n4313_o;
  wire n4314_o;
  wire n4315_o;
  wire n4316_o;
  wire n4318_o;
  wire n4319_o;
  wire n4320_o;
  wire n4321_o;
  wire n4323_o;
  wire n4324_o;
  wire n4325_o;
  wire n4326_o;
  wire n4328_o;
  wire n4329_o;
  wire n4330_o;
  wire n4331_o;
  wire n4333_o;
  wire n4334_o;
  wire n4335_o;
  wire n4336_o;
  wire n4338_o;
  wire n4339_o;
  wire n4340_o;
  wire n4341_o;
  wire n4343_o;
  wire n4344_o;
  wire n4345_o;
  wire n4346_o;
  wire n4348_o;
  wire n4349_o;
  wire n4350_o;
  wire n4351_o;
  wire n4353_o;
  wire n4354_o;
  wire n4355_o;
  wire n4356_o;
  wire n4358_o;
  wire n4359_o;
  wire n4360_o;
  wire n4361_o;
  wire n4363_o;
  wire n4364_o;
  wire n4365_o;
  wire n4366_o;
  wire n4368_o;
  wire n4369_o;
  wire n4370_o;
  wire n4371_o;
  wire n4373_o;
  wire n4374_o;
  wire n4375_o;
  wire n4376_o;
  wire n4378_o;
  wire n4379_o;
  wire n4380_o;
  wire n4381_o;
  wire n4383_o;
  wire n4384_o;
  wire n4385_o;
  wire n4386_o;
  wire n4388_o;
  wire n4389_o;
  wire n4390_o;
  wire n4391_o;
  wire n4393_o;
  wire n4394_o;
  wire n4395_o;
  wire n4396_o;
  wire n4398_o;
  wire n4399_o;
  wire n4400_o;
  wire n4401_o;
  wire n4403_o;
  wire n4404_o;
  wire n4405_o;
  wire n4406_o;
  wire n4408_o;
  wire n4409_o;
  wire n4410_o;
  wire n4411_o;
  wire n4413_o;
  wire n4414_o;
  wire n4415_o;
  wire n4416_o;
  wire n4418_o;
  wire n4419_o;
  wire n4420_o;
  wire n4421_o;
  wire n4423_o;
  wire n4424_o;
  wire n4425_o;
  wire n4426_o;
  wire n4428_o;
  wire n4429_o;
  wire n4430_o;
  wire n4431_o;
  wire n4433_o;
  wire n4434_o;
  wire n4435_o;
  wire n4438_o;
  wire n4439_o;
  wire n4440_o;
  wire n4441_o;
  wire n4442_o;
  wire n4443_o;
  wire n4444_o;
  wire n4445_o;
  wire n4446_o;
  wire n4447_o;
  wire n4448_o;
  wire n4449_o;
  wire n4450_o;
  wire n4451_o;
  wire n4452_o;
  wire n4453_o;
  wire n4454_o;
  wire n4455_o;
  wire n4456_o;
  wire n4457_o;
  wire n4458_o;
  wire n4459_o;
  wire n4460_o;
  wire n4461_o;
  wire n4462_o;
  wire n4463_o;
  wire n4464_o;
  wire n4465_o;
  wire n4466_o;
  wire n4467_o;
  wire n4468_o;
  wire n4469_o;
  wire n4470_o;
  wire n4471_o;
  wire n4472_o;
  wire n4473_o;
  wire n4474_o;
  wire n4475_o;
  wire n4476_o;
  wire n4477_o;
  wire n4478_o;
  wire n4479_o;
  wire n4480_o;
  wire n4481_o;
  wire n4482_o;
  wire n4483_o;
  wire n4484_o;
  wire n4485_o;
  wire n4486_o;
  wire n4487_o;
  wire n4488_o;
  wire n4489_o;
  wire n4490_o;
  wire n4491_o;
  wire n4492_o;
  wire n4493_o;
  wire n4494_o;
  wire n4495_o;
  wire n4496_o;
  wire n4497_o;
  wire n4498_o;
  wire n4499_o;
  wire n4500_o;
  wire n4501_o;
  wire n4502_o;
  wire n4503_o;
  wire n4504_o;
  wire n4505_o;
  wire n4506_o;
  wire n4507_o;
  wire n4508_o;
  wire n4509_o;
  wire n4510_o;
  wire n4511_o;
  wire n4512_o;
  wire n4513_o;
  wire n4514_o;
  wire n4515_o;
  wire n4516_o;
  wire n4517_o;
  wire n4518_o;
  wire n4519_o;
  wire n4520_o;
  wire n4521_o;
  wire n4522_o;
  wire n4523_o;
  wire n4524_o;
  wire n4525_o;
  wire n4526_o;
  wire n4527_o;
  wire n4528_o;
  wire n4529_o;
  wire n4530_o;
  wire n4531_o;
  wire n4532_o;
  wire n4533_o;
  wire n4534_o;
  wire n4535_o;
  wire n4536_o;
  wire n4537_o;
  wire n4538_o;
  wire n4539_o;
  wire n4540_o;
  wire n4541_o;
  wire n4542_o;
  wire n4543_o;
  wire n4544_o;
  wire n4545_o;
  wire n4546_o;
  wire n4547_o;
  wire n4548_o;
  wire n4549_o;
  wire n4550_o;
  wire n4551_o;
  wire n4552_o;
  wire n4553_o;
  wire n4554_o;
  wire n4555_o;
  wire n4556_o;
  wire n4557_o;
  wire n4558_o;
  wire n4559_o;
  wire n4560_o;
  wire n4561_o;
  wire n4562_o;
  wire n4563_o;
  wire n4564_o;
  wire n4565_o;
  wire n4566_o;
  wire n4567_o;
  wire n4568_o;
  wire n4569_o;
  wire n4570_o;
  wire [41:0] n4573_o;
  wire [41:0] n4576_o;
  wire n4580_o;
  wire n4583_o;
  wire n4585_o;
  wire n4587_o;
  wire n4589_o;
  wire n4590_o;
  wire [5:0] n4592_o;
  wire n4593_o;
  wire [6:0] n4594_o;
  wire n4595_o;
  wire n4597_o;
  wire n4599_o;
  wire n4601_o;
  wire n4603_o;
  wire n4605_o;
  wire n4607_o;
  wire n4609_o;
  wire n4611_o;
  wire n4613_o;
  wire n4615_o;
  wire n4617_o;
  wire n4619_o;
  wire n4621_o;
  wire n4623_o;
  wire n4625_o;
  wire n4627_o;
  wire n4629_o;
  wire n4631_o;
  wire n4633_o;
  wire n4635_o;
  wire n4637_o;
  wire n4639_o;
  wire n4641_o;
  wire n4643_o;
  wire n4645_o;
  wire n4647_o;
  wire [6:0] n4651_o;
  wire [6:0] n4652_o;
  wire [6:0] n4653_o;
  wire [6:0] n4654_o;
  wire [6:0] n4655_o;
  wire [6:0] n4656_o;
  wire [6:0] n4657_o;
  wire [6:0] n4658_o;
  wire [6:0] n4659_o;
  wire [6:0] n4660_o;
  wire [6:0] n4661_o;
  wire [6:0] n4662_o;
  wire [6:0] n4663_o;
  wire [6:0] n4664_o;
  wire [6:0] n4665_o;
  wire [6:0] n4666_o;
  wire [6:0] n4667_o;
  wire [6:0] n4668_o;
  wire [6:0] n4669_o;
  wire [6:0] n4670_o;
  wire [6:0] n4671_o;
  wire [6:0] n4672_o;
  wire [6:0] n4673_o;
  wire [6:0] n4674_o;
  wire [6:0] n4675_o;
  wire [6:0] n4676_o;
  wire [6:0] n4677_o;
  wire [6:0] n4678_o;
  wire [6:0] n4679_o;
  wire [6:0] n4680_o;
  wire [6:0] n4681_o;
  wire n4687_o;
  wire n4690_o;
  wire n4691_o;
  wire n4692_o;
  wire n4693_o;
  wire [3:0] n4694_o;
  wire n4696_o;
  wire n4697_o;
  wire n4698_o;
  wire n4700_o;
  wire n4701_o;
  wire n4702_o;
  wire n4704_o;
  wire n4705_o;
  wire n4706_o;
  wire n4718_o;
  wire n4720_o;
  wire n4722_o;
  wire n4723_o;
  wire n4724_o;
  wire n4725_o;
  wire n4726_o;
  wire n4727_o;
  wire n4728_o;
  wire n4729_o;
  wire n4730_o;
  wire n4731_o;
  wire n4732_o;
  wire n4733_o;
  wire n4734_o;
  wire n4735_o;
  wire n4736_o;
  wire n4737_o;
  wire n4738_o;
  wire n4739_o;
  wire n4740_o;
  wire n4741_o;
  wire n4742_o;
  wire n4743_o;
  wire n4744_o;
  wire n4745_o;
  wire n4746_o;
  wire n4747_o;
  wire n4748_o;
  wire n4749_o;
  wire n4750_o;
  wire n4751_o;
  wire n4752_o;
  wire n4753_o;
  wire n4754_o;
  wire n4755_o;
  wire n4756_o;
  wire n4757_o;
  wire n4758_o;
  wire n4759_o;
  wire n4760_o;
  wire n4761_o;
  wire n4762_o;
  wire n4763_o;
  wire n4764_o;
  wire n4765_o;
  wire n4774_o;
  wire n4776_o;
  wire n4778_o;
  wire n4779_o;
  wire n4780_o;
  wire n4781_o;
  wire n4782_o;
  wire n4783_o;
  wire n4784_o;
  wire n4785_o;
  wire n4786_o;
  wire n4787_o;
  wire n4788_o;
  wire n4789_o;
  wire n4790_o;
  wire n4791_o;
  wire n4792_o;
  wire n4793_o;
  wire n4794_o;
  wire n4795_o;
  wire n4796_o;
  wire n4797_o;
  wire n4798_o;
  wire n4808_o;
  wire n4810_o;
  wire n4812_o;
  wire n4813_o;
  wire n4814_o;
  wire n4815_o;
  wire n4816_o;
  wire n4817_o;
  wire n4818_o;
  wire n4819_o;
  wire n4820_o;
  wire n4821_o;
  wire n4822_o;
  wire n4823_o;
  wire n4824_o;
  wire n4825_o;
  wire n4826_o;
  wire n4827_o;
  wire n4828_o;
  wire n4829_o;
  wire n4830_o;
  wire n4831_o;
  wire n4832_o;
  wire n4833_o;
  wire n4834_o;
  wire n4835_o;
  wire n4836_o;
  wire n4837_o;
  wire n4838_o;
  wire n4839_o;
  wire n4840_o;
  wire n4841_o;
  wire n4842_o;
  wire n4843_o;
  wire n4844_o;
  wire n4845_o;
  wire n4846_o;
  wire n4847_o;
  wire n4848_o;
  wire n4849_o;
  wire n4850_o;
  wire n4851_o;
  wire n4852_o;
  wire n4853_o;
  wire n4854_o;
  wire n4855_o;
  wire n4856_o;
  wire n4857_o;
  wire n4858_o;
  wire n4859_o;
  wire n4860_o;
  wire n4861_o;
  wire n4862_o;
  wire n4863_o;
  wire [31:0] n4865_o;
  wire n4866_o;
  wire [31:0] n4867_o;
  wire [31:0] n4868_o;
  wire [11:0] n4869_o;
  wire [1:0] n4870_o;
  wire n4871_o;
  wire [2:0] n4872_o;
  wire n4873_o;
  wire [3:0] n4874_o;
  wire [7:0] n4875_o;
  wire [11:0] n4876_o;
  wire [2:0] n4877_o;
  wire n4880_o;
  wire [4:0] n4881_o;
  localparam [31:0] n4882_o = 32'b00000000000000000000000000000000;
  wire [26:0] n4883_o;
  wire [31:0] n4884_o;
  wire [31:0] n4885_o;
  wire [1:0] n4886_o;
  wire n4888_o;
  wire [31:0] n4889_o;
  wire [31:0] n4890_o;
  wire [1:0] n4892_o;
  wire [31:0] n4893_o;
  wire [31:0] n4894_o;
  wire [31:0] n4895_o;
  wire n4897_o;
  wire [31:0] n4898_o;
  wire [31:0] n4899_o;
  wire [31:0] n4900_o;
  wire n4902_o;
  wire [31:0] n4903_o;
  wire [1:0] n4904_o;
  reg [31:0] n4905_o;
  wire n4906_o;
  wire [11:0] n4907_o;
  wire [31:0] n4908_o;
  wire n4910_o;
  wire n4942_o;
  wire n4943_o;
  wire n4944_o;
  wire n4945_o;
  wire n4946_o;
  wire [11:0] n4947_o;
  wire n4948_o;
  wire n4949_o;
  wire n4950_o;
  wire n4951_o;
  wire n4952_o;
  wire n4953_o;
  wire n4954_o;
  wire n4956_o;
  wire n4957_o;
  wire n4958_o;
  wire n4959_o;
  wire [15:0] n4960_o;
  wire n4962_o;
  wire [1:0] n4963_o;
  wire n4965_o;
  wire [24:0] n4966_o;
  wire [29:0] n4968_o;
  wire [31:0] n4970_o;
  wire [29:0] n4971_o;
  wire [31:0] n4973_o;
  wire [31:0] n4974_o;
  wire n4976_o;
  wire n4977_o;
  wire n4978_o;
  wire n4979_o;
  wire n4981_o;
  wire [31:0] n4982_o;
  wire n4984_o;
  wire [30:0] n4985_o;
  wire [31:0] n4987_o;
  wire n4989_o;
  wire n4990_o;
  wire [4:0] n4991_o;
  wire [5:0] n4992_o;
  wire n4994_o;
  wire n4995_o;
  wire n4996_o;
  wire n4998_o;
  wire n5000_o;
  wire n5002_o;
  wire n5004_o;
  wire n5006_o;
  wire n5008_o;
  wire [12:0] n5009_o;
  wire n5010_o;
  reg n5011_o;
  wire n5012_o;
  reg n5013_o;
  wire n5014_o;
  reg n5015_o;
  wire n5016_o;
  reg n5017_o;
  wire n5018_o;
  reg n5019_o;
  wire n5020_o;
  reg n5021_o;
  wire n5022_o;
  reg n5023_o;
  wire n5024_o;
  reg n5025_o;
  wire [15:0] n5026_o;
  reg [15:0] n5027_o;
  wire [31:0] n5028_o;
  reg [31:0] n5029_o;
  wire [5:0] n5030_o;
  reg [5:0] n5031_o;
  wire [31:0] n5032_o;
  reg [31:0] n5033_o;
  wire [31:0] n5034_o;
  reg [31:0] n5035_o;
  wire n5036_o;
  reg n5037_o;
  wire n5038_o;
  reg n5039_o;
  wire n5040_o;
  reg n5041_o;
  wire n5042_o;
  wire n5043_o;
  wire [4:0] n5044_o;
  wire [5:0] n5045_o;
  wire [30:0] n5046_o;
  wire [31:0] n5048_o;
  wire n5049_o;
  wire n5050_o;
  wire n5051_o;
  wire n5052_o;
  wire [31:0] n5054_o;
  wire n5055_o;
  wire n5056_o;
  wire n5058_o;
  wire n5060_o;
  wire n5062_o;
  wire n5063_o;
  wire [29:0] n5064_o;
  wire n5065_o;
  wire [31:0] n5067_o;
  wire [31:0] n5068_o;
  wire n5071_o;
  wire n5072_o;
  wire n5073_o;
  wire n5074_o;
  wire n5076_o;
  wire n5078_o;
  wire n5080_o;
  wire n5081_o;
  wire n5082_o;
  wire [3:0] n5084_o;
  wire [3:0] n5085_o;
  wire [3:0] n5086_o;
  wire n5087_o;
  wire n5088_o;
  wire [2:0] n5089_o;
  wire [37:0] n5090_o;
  wire [63:0] n5091_o;
  wire [2:0] n5092_o;
  wire [2:0] n5093_o;
  wire n5094_o;
  wire n5095_o;
  wire n5096_o;
  wire n5097_o;
  wire [37:0] n5098_o;
  wire [37:0] n5099_o;
  wire [63:0] n5100_o;
  wire [63:0] n5101_o;
  wire [3:0] n5102_o;
  wire [23:0] n5103_o;
  wire [69:0] n5104_o;
  wire [33:0] n5105_o;
  wire [3:0] n5106_o;
  wire [3:0] n5107_o;
  wire [19:0] n5108_o;
  wire [19:0] n5109_o;
  wire [19:0] n5110_o;
  wire n5111_o;
  wire n5112_o;
  wire [37:0] n5113_o;
  wire [37:0] n5114_o;
  wire [31:0] n5115_o;
  wire [31:0] n5116_o;
  wire [31:0] n5117_o;
  wire [63:0] n5118_o;
  wire [63:0] n5119_o;
  wire [33:0] n5120_o;
  wire [33:0] n5121_o;
  wire n5122_o;
  wire n5123_o;
  wire [23:0] n5137_o;
  wire [189:0] n5138_o;
  wire [63:0] n5139_o;
  wire [2:0] n5140_o;
  wire [23:0] n5155_o;
  wire [189:0] n5156_o;
  wire [63:0] n5157_o;
  wire [2:0] n5158_o;
  wire n5168_o;
  wire n5169_o;
  wire n5170_o;
  wire [11:0] n5171_o;
  wire n5173_o;
  wire n5174_o;
  wire n5175_o;
  wire n5178_o;
  wire n5179_o;
  wire n5180_o;
  wire [11:0] n5181_o;
  wire n5183_o;
  wire n5184_o;
  wire n5185_o;
  wire n5188_o;
  wire n5189_o;
  wire n5190_o;
  wire [11:0] n5192_o;
  wire n5193_o;
  wire n5194_o;
  wire n5195_o;
  wire n5196_o;
  wire [1:0] n5197_o;
  wire n5198_o;
  wire n5199_o;
  wire n5202_o;
  wire n5204_o;
  localparam [1:0] n5220_o = 2'b01;
  wire n5222_o;
  wire n5223_o;
  wire n5224_o;
  wire n5225_o;
  wire [15:0] n5226_o;
  wire n5228_o;
  wire [31:0] n5229_o;
  wire n5231_o;
  wire n5232_o;
  wire n5233_o;
  wire n5235_o;
  wire [31:0] n5236_o;
  wire n5238_o;
  wire [30:0] n5239_o;
  wire [31:0] n5241_o;
  wire n5243_o;
  wire n5244_o;
  wire [4:0] n5245_o;
  wire n5247_o;
  wire [31:0] n5248_o;
  wire n5250_o;
  wire n5251_o;
  wire n5252_o;
  wire n5253_o;
  wire [15:0] n5254_o;
  wire n5256_o;
  wire [31:0] n5257_o;
  wire n5259_o;
  wire n5260_o;
  wire n5261_o;
  wire n5263_o;
  wire n5265_o;
  wire n5267_o;
  wire n5269_o;
  wire n5271_o;
  wire n5273_o;
  wire n5275_o;
  wire n5277_o;
  wire n5279_o;
  wire n5281_o;
  wire n5283_o;
  wire n5285_o;
  wire n5287_o;
  wire n5289_o;
  wire [31:0] n5290_o;
  wire n5292_o;
  wire n5294_o;
  wire n5295_o;
  wire [31:0] n5296_o;
  wire n5298_o;
  wire n5300_o;
  wire n5301_o;
  wire n5303_o;
  wire n5305_o;
  wire n5306_o;
  wire n5308_o;
  wire n5310_o;
  wire n5311_o;
  wire n5313_o;
  wire n5315_o;
  wire n5316_o;
  wire n5318_o;
  wire n5320_o;
  wire n5321_o;
  wire n5323_o;
  wire n5325_o;
  wire n5326_o;
  wire n5328_o;
  wire n5330_o;
  wire n5331_o;
  wire n5333_o;
  wire n5335_o;
  wire n5336_o;
  wire n5338_o;
  wire n5340_o;
  wire n5341_o;
  wire n5343_o;
  wire n5345_o;
  wire n5346_o;
  wire n5348_o;
  wire n5350_o;
  wire n5351_o;
  wire n5353_o;
  wire n5355_o;
  wire n5356_o;
  wire n5358_o;
  wire n5360_o;
  wire n5361_o;
  wire n5363_o;
  wire n5365_o;
  wire n5366_o;
  wire [31:0] n5367_o;
  wire n5369_o;
  wire n5371_o;
  wire n5372_o;
  wire [31:0] n5373_o;
  wire n5375_o;
  wire n5377_o;
  wire n5378_o;
  wire n5380_o;
  wire n5382_o;
  wire n5383_o;
  wire n5385_o;
  wire n5387_o;
  wire n5388_o;
  wire n5390_o;
  wire n5392_o;
  wire n5393_o;
  wire n5395_o;
  wire n5397_o;
  wire n5398_o;
  wire n5400_o;
  wire n5402_o;
  wire n5403_o;
  wire n5405_o;
  wire n5407_o;
  wire n5408_o;
  wire n5410_o;
  wire n5412_o;
  wire n5413_o;
  wire n5415_o;
  wire n5417_o;
  wire n5418_o;
  wire n5420_o;
  wire n5422_o;
  wire n5423_o;
  wire n5425_o;
  wire n5427_o;
  wire n5428_o;
  wire n5430_o;
  wire n5432_o;
  wire n5433_o;
  wire n5435_o;
  wire n5437_o;
  wire n5438_o;
  wire n5440_o;
  wire n5442_o;
  wire n5443_o;
  wire n5445_o;
  localparam [4:0] n5446_o = 5'b10011;
  wire n5448_o;
  wire n5450_o;
  wire n5452_o;
  wire n5454_o;
  wire n5456_o;
  wire n5458_o;
  wire n5460_o;
  wire n5462_o;
  wire n5464_o;
  wire n5495_o;
  wire [65:0] n5496_o;
  wire n5497_o;
  wire n5498_o;
  wire n5499_o;
  wire n5500_o;
  wire n5501_o;
  wire n5502_o;
  wire n5503_o;
  wire n5504_o;
  wire n5505_o;
  wire n5506_o;
  wire n5508_o;
  reg n5512_o;
  wire n5513_o;
  wire n5514_o;
  wire n5515_o;
  wire n5516_o;
  wire n5517_o;
  wire n5518_o;
  wire n5519_o;
  wire n5520_o;
  wire n5521_o;
  wire n5522_o;
  wire n5524_o;
  reg n5528_o;
  wire n5529_o;
  wire n5530_o;
  wire n5531_o;
  wire n5532_o;
  wire n5533_o;
  wire n5534_o;
  wire n5535_o;
  wire n5536_o;
  wire n5537_o;
  wire n5538_o;
  wire n5540_o;
  reg n5544_o;
  wire n5545_o;
  wire n5546_o;
  wire n5547_o;
  wire n5548_o;
  wire n5549_o;
  wire n5550_o;
  wire n5551_o;
  wire n5552_o;
  wire n5553_o;
  wire n5554_o;
  wire n5556_o;
  reg n5560_o;
  wire n5561_o;
  wire n5562_o;
  wire n5563_o;
  wire n5564_o;
  wire n5565_o;
  wire n5566_o;
  wire n5567_o;
  wire n5568_o;
  wire n5569_o;
  wire n5570_o;
  wire n5572_o;
  reg n5576_o;
  wire n5577_o;
  wire n5578_o;
  wire n5579_o;
  wire n5580_o;
  wire n5581_o;
  wire n5582_o;
  wire n5583_o;
  wire n5584_o;
  wire n5585_o;
  reg n5590_o;
  wire n5591_o;
  wire n5592_o;
  wire n5593_o;
  wire n5594_o;
  wire n5595_o;
  wire n5596_o;
  wire n5597_o;
  wire n5598_o;
  wire n5599_o;
  reg n5604_o;
  wire n5605_o;
  wire n5606_o;
  wire n5607_o;
  wire n5608_o;
  wire n5609_o;
  wire n5610_o;
  wire n5611_o;
  wire n5612_o;
  wire n5613_o;
  reg n5618_o;
  wire n5619_o;
  wire n5620_o;
  wire n5621_o;
  wire n5622_o;
  wire n5623_o;
  wire n5624_o;
  wire n5625_o;
  wire n5626_o;
  wire n5627_o;
  reg n5632_o;
  wire n5633_o;
  wire n5634_o;
  wire n5635_o;
  wire n5636_o;
  wire n5637_o;
  wire n5638_o;
  wire n5639_o;
  wire n5640_o;
  wire n5641_o;
  reg n5646_o;
  wire n5647_o;
  wire n5648_o;
  wire n5649_o;
  wire n5650_o;
  wire n5651_o;
  wire n5652_o;
  wire n5653_o;
  wire n5654_o;
  wire n5655_o;
  reg n5660_o;
  wire n5661_o;
  wire n5662_o;
  wire n5663_o;
  wire n5664_o;
  wire n5665_o;
  wire n5666_o;
  wire n5667_o;
  wire n5668_o;
  wire n5669_o;
  wire n5670_o;
  reg n5675_o;
  wire n5676_o;
  wire n5677_o;
  wire n5678_o;
  wire n5679_o;
  wire n5680_o;
  wire n5681_o;
  wire n5682_o;
  wire n5683_o;
  wire n5684_o;
  wire n5685_o;
  reg n5690_o;
  wire [2:0] n5691_o;
  wire [2:0] n5692_o;
  wire [2:0] n5693_o;
  wire [2:0] n5694_o;
  wire [2:0] n5695_o;
  wire [2:0] n5696_o;
  wire [2:0] n5697_o;
  wire [2:0] n5698_o;
  wire [2:0] n5699_o;
  reg [2:0] n5704_o;
  wire n5705_o;
  wire n5706_o;
  wire n5707_o;
  wire n5708_o;
  wire n5709_o;
  wire n5710_o;
  wire n5711_o;
  wire n5712_o;
  wire n5713_o;
  wire n5714_o;
  wire n5715_o;
  reg n5720_o;
  wire n5721_o;
  wire n5722_o;
  wire n5723_o;
  wire n5724_o;
  wire n5725_o;
  wire n5726_o;
  wire n5727_o;
  wire n5728_o;
  wire n5729_o;
  wire n5730_o;
  wire n5731_o;
  reg n5736_o;
  wire [1:0] n5737_o;
  wire [1:0] n5738_o;
  wire [1:0] n5739_o;
  wire [1:0] n5740_o;
  wire [1:0] n5741_o;
  wire [1:0] n5742_o;
  wire [1:0] n5743_o;
  wire [1:0] n5744_o;
  wire [1:0] n5745_o;
  wire [1:0] n5746_o;
  wire [1:0] n5747_o;
  reg [1:0] n5752_o;
  wire n5753_o;
  wire n5754_o;
  wire n5755_o;
  wire n5756_o;
  wire n5757_o;
  wire n5758_o;
  wire n5759_o;
  wire n5760_o;
  wire n5761_o;
  wire n5762_o;
  wire n5763_o;
  reg n5768_o;
  wire n5769_o;
  wire n5770_o;
  wire n5771_o;
  wire n5772_o;
  wire n5773_o;
  wire n5774_o;
  wire n5775_o;
  wire n5776_o;
  wire n5777_o;
  wire n5778_o;
  wire n5779_o;
  reg n5784_o;
  wire n5785_o;
  wire n5786_o;
  wire n5787_o;
  wire n5788_o;
  wire n5789_o;
  wire n5790_o;
  wire n5791_o;
  wire n5792_o;
  wire n5793_o;
  wire n5794_o;
  wire n5795_o;
  reg n5800_o;
  wire n5801_o;
  wire n5802_o;
  wire n5803_o;
  wire n5804_o;
  wire n5805_o;
  wire n5806_o;
  wire n5807_o;
  wire n5808_o;
  wire n5809_o;
  wire n5810_o;
  wire n5811_o;
  reg n5816_o;
  wire [4:0] n5817_o;
  wire [4:0] n5818_o;
  wire [4:0] n5819_o;
  wire [4:0] n5820_o;
  wire [4:0] n5821_o;
  wire [4:0] n5822_o;
  wire [4:0] n5823_o;
  wire [4:0] n5824_o;
  wire [4:0] n5825_o;
  wire [4:0] n5826_o;
  wire [4:0] n5827_o;
  reg [4:0] n5832_o;
  wire n5833_o;
  wire n5834_o;
  wire n5835_o;
  wire n5836_o;
  wire n5837_o;
  wire n5838_o;
  wire n5839_o;
  wire n5840_o;
  wire n5841_o;
  wire n5842_o;
  wire n5843_o;
  reg n5848_o;
  wire n5849_o;
  wire n5850_o;
  wire n5851_o;
  wire n5852_o;
  wire n5853_o;
  wire n5854_o;
  wire n5855_o;
  wire n5856_o;
  wire n5857_o;
  wire n5858_o;
  wire n5859_o;
  wire n5860_o;
  reg n5865_o;
  wire n5866_o;
  wire n5867_o;
  wire n5868_o;
  wire n5869_o;
  wire n5870_o;
  wire n5871_o;
  wire n5872_o;
  wire n5873_o;
  wire n5874_o;
  wire n5875_o;
  wire n5876_o;
  wire n5877_o;
  reg n5882_o;
  wire n5910_o;
  wire n5914_o;
  wire n5915_o;
  wire [31:0] n5916_o;
  wire [31:0] n5918_o;
  wire [31:0] n5926_o;
  localparam [15:0] n5928_o = 16'b0000000000000000;
  localparam [15:0] n5929_o = 16'b0000000000000000;
  wire n5930_o;
  wire [3:0] n5931_o;
  wire n5933_o;
  wire n5934_o;
  wire n5935_o;
  wire n5936_o;
  wire [3:0] n5937_o;
  wire [3:0] n5942_o;
  wire [15:0] n5947_o;
  wire [15:0] n5948_o;
  wire [31:0] n5949_o;
  wire [31:0] n5950_o;
  wire [31:0] n5951_o;
  wire n5954_o;
  wire n5959_o;
  wire [31:0] n5960_o;
  wire [31:0] n5961_o;
  wire [31:0] n5962_o;
  wire n5963_o;
  wire n5964_o;
  wire [31:0] n5965_o;
  wire [31:0] n5966_o;
  wire n5967_o;
  wire [31:0] n5968_o;
  wire [31:0] n5969_o;
  wire [31:0] n5970_o;
  wire [31:0] n5981_o;
  wire [32:0] n5983_o;
  wire [32:0] n5985_o;
  wire n5986_o;
  wire [32:0] n5987_o;
  wire [31:0] n5988_o;
  wire [32:0] n5990_o;
  wire [32:0] n5992_o;
  wire n5994_o;
  wire n5999_o;
  wire [31:0] n6000_o;
  wire [31:0] n6001_o;
  wire [31:0] n6002_o;
  wire n6003_o;
  wire n6004_o;
  wire [31:0] n6005_o;
  wire [31:0] n6006_o;
  wire n6007_o;
  wire [31:0] n6008_o;
  wire [31:0] n6009_o;
  wire [31:0] n6010_o;
  wire [31:0] n6021_o;
  wire [32:0] n6023_o;
  wire [32:0] n6025_o;
  wire n6026_o;
  wire [32:0] n6027_o;
  wire [31:0] n6028_o;
  wire [32:0] n6030_o;
  wire [32:0] n6032_o;
  wire n6034_o;
  wire n6039_o;
  wire [31:0] n6040_o;
  wire [31:0] n6041_o;
  wire [31:0] n6042_o;
  wire n6043_o;
  wire n6044_o;
  wire [31:0] n6045_o;
  wire [31:0] n6046_o;
  wire n6047_o;
  wire [31:0] n6048_o;
  wire [31:0] n6049_o;
  wire [31:0] n6050_o;
  wire [31:0] n6061_o;
  wire [32:0] n6063_o;
  wire [32:0] n6065_o;
  wire n6066_o;
  wire [32:0] n6067_o;
  wire [31:0] n6068_o;
  wire [32:0] n6070_o;
  wire [32:0] n6072_o;
  wire [31:0] n6074_o;
  localparam [95:0] n6075_o = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n6077_o;
  localparam [95:0] n6078_o = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n6080_o;
  wire [31:0] n6081_o;
  wire [31:0] n6082_o;
  wire [31:0] n6083_o;
  wire n6088_o;
  localparam [15:0] n6091_o = 16'b0000000000000000;
  wire n6092_o;
  wire n6093_o;
  wire n6094_o;
  wire n6095_o;
  wire n6096_o;
  wire n6097_o;
  wire n6098_o;
  wire n6100_o;
  wire n6101_o;
  wire n6102_o;
  wire n6103_o;
  wire n6104_o;
  wire n6105_o;
  wire n6106_o;
  wire [12:0] n6107_o;
  wire n6108_o;
  wire [15:0] n6109_o;
  wire n6115_o;
  wire n6116_o;
  wire [3:0] n6120_o;
  wire n6122_o;
  wire n6123_o;
  wire [3:0] n6126_o;
  wire n6128_o;
  wire n6129_o;
  wire n6130_o;
  wire n6131_o;
  wire [3:0] n6134_o;
  wire n6136_o;
  wire [1:0] n6137_o;
  wire n6139_o;
  wire n6140_o;
  wire n6141_o;
  wire [3:0] n6144_o;
  wire n6146_o;
  wire n6147_o;
  wire [3:0] n6150_o;
  wire n6152_o;
  wire n6153_o;
  wire [3:0] n6156_o;
  wire n6158_o;
  wire n6159_o;
  wire n6162_o;
  wire n6163_o;
  wire n6164_o;
  wire n6165_o;
  wire n6166_o;
  wire n6169_o;
  wire n6170_o;
  wire n6171_o;
  wire n6172_o;
  wire n6175_o;
  wire n6176_o;
  wire [3:0] n6177_o;
  wire n6179_o;
  wire n6180_o;
  wire n6181_o;
  wire n6184_o;
  wire n6185_o;
  wire n6194_o;
  wire n6197_o;
  wire n6199_o;
  wire [2:0] n6204_o;
  wire n6208_o;
  wire n6209_o;
  wire n6210_o;
  wire [1:0] n6211_o;
  wire n6215_o;
  wire n6223_o;
  wire [3:0] n6225_o;
  wire n6233_o;
  reg n6236_q;
  reg [34:0] n6237_q;
  wire [37:0] n6238_o;
  wire [75:0] n6239_o;
  reg n6240_q;
  wire [87:0] n6241_o;
  wire [16:0] n6242_o;
  wire [31:0] n6243_o;
  wire [31:0] n6244_o;
  reg [31:0] n6245_q;
  reg [31:0] n6246_q;
  wire [31:0] n6247_o;
  wire [31:0] n6248_o;
  reg [31:0] n6249_q;
  reg n6250_q;
  reg [31:0] n6251_q;
  reg [3:0] n6252_q;
  wire [203:0] n6253_o;
  reg [9:0] n6254_q;
  wire [20:0] n6255_o;
  reg n6256_q;
  reg n6257_q;
  reg [6:0] n6258_q;
  reg [41:0] n6259_q;
  reg [10:0] n6260_q;
  wire [103:0] n6261_o;
  reg [66:0] n6262_q;
  wire [66:0] n6263_o;
  reg [31:0] n6264_q;
  reg n6265_q;
  reg [31:0] n6266_q;
  reg [2:0] n6267_q;
  reg [63:0] n6268_q;
  reg [189:0] n6269_q;
  reg n6270_q;
  reg [23:0] n6271_q;
  reg n6272_q;
  wire [507:0] n6273_o;
  reg [15:0] n6275_q;
  reg n6276_q;
  reg [31:0] n6277_q;
  reg [31:0] n6278_q;
  reg n6279_q;
  reg [31:0] n6280_q;
  reg [31:0] n6281_q;
  reg n6282_q;
  reg [31:0] n6283_q;
  reg [31:0] n6284_q;
  wire [341:0] n6285_o;
  wire [95:0] n6286_o;
  wire [95:0] n6287_o;
  wire [11:0] n6288_o;
  wire [4:0] n6289_o;
  wire [31:0] n6290_o;
  wire [66:0] n6291_o;
  wire [73:0] n6292_o;
  reg [31:0] n6293_q;
  wire n6294_o;
  wire n6295_o;
  wire n6296_o;
  wire n6297_o;
  wire n6298_o;
  wire n6299_o;
  wire n6300_o;
  wire n6301_o;
  wire n6302_o;
  wire n6303_o;
  wire n6304_o;
  wire n6305_o;
  wire n6306_o;
  wire n6307_o;
  wire n6308_o;
  wire n6309_o;
  wire n6310_o;
  wire n6311_o;
  wire n6312_o;
  wire n6313_o;
  wire n6314_o;
  wire n6315_o;
  wire n6316_o;
  wire n6317_o;
  wire n6318_o;
  wire n6319_o;
  wire n6320_o;
  wire n6321_o;
  wire n6322_o;
  wire n6323_o;
  wire n6324_o;
  wire n6325_o;
  wire n6326_o;
  wire n6327_o;
  wire n6328_o;
  wire n6329_o;
  wire n6330_o;
  wire n6331_o;
  wire n6332_o;
  wire n6333_o;
  wire n6334_o;
  wire n6335_o;
  wire n6336_o;
  wire n6337_o;
  wire n6338_o;
  wire n6339_o;
  wire n6340_o;
  wire n6341_o;
  wire n6342_o;
  wire n6343_o;
  wire n6344_o;
  wire n6345_o;
  wire n6346_o;
  wire n6347_o;
  wire n6348_o;
  wire n6349_o;
  wire n6350_o;
  wire n6351_o;
  wire n6352_o;
  wire n6353_o;
  wire n6354_o;
  wire n6355_o;
  wire n6356_o;
  wire n6357_o;
  wire n6358_o;
  wire n6359_o;
  wire n6360_o;
  wire n6361_o;
  wire [15:0] n6362_o;
  wire n6363_o;
  wire n6364_o;
  wire n6365_o;
  wire n6366_o;
  wire n6367_o;
  wire n6368_o;
  wire n6369_o;
  wire n6370_o;
  wire n6371_o;
  wire n6372_o;
  wire n6373_o;
  wire n6374_o;
  wire n6375_o;
  wire n6376_o;
  wire n6377_o;
  wire n6378_o;
  wire n6379_o;
  wire n6380_o;
  wire n6381_o;
  wire n6382_o;
  wire n6383_o;
  wire n6384_o;
  wire n6385_o;
  wire n6386_o;
  wire n6387_o;
  wire n6388_o;
  wire n6389_o;
  wire n6390_o;
  wire n6391_o;
  wire n6392_o;
  wire n6393_o;
  wire n6394_o;
  wire n6395_o;
  wire n6396_o;
  wire n6397_o;
  wire n6398_o;
  wire n6399_o;
  wire n6400_o;
  wire n6401_o;
  wire n6402_o;
  wire n6403_o;
  wire n6404_o;
  wire n6405_o;
  wire n6406_o;
  wire n6407_o;
  wire n6408_o;
  wire n6409_o;
  wire n6410_o;
  wire n6411_o;
  wire n6412_o;
  wire n6413_o;
  wire n6414_o;
  wire n6415_o;
  wire n6416_o;
  wire n6417_o;
  wire n6418_o;
  wire n6419_o;
  wire n6420_o;
  wire n6421_o;
  wire n6422_o;
  wire n6423_o;
  wire n6424_o;
  wire n6425_o;
  wire n6426_o;
  wire n6427_o;
  wire n6428_o;
  wire n6429_o;
  wire n6430_o;
  wire [15:0] n6431_o;
  assign ctrl_o_rf_wb_en = n2328_o; //(module output)
  assign ctrl_o_rf_rs1 = n2329_o; //(module output)
  assign ctrl_o_rf_rs2 = n2330_o; //(module output)
  assign ctrl_o_rf_rs3 = n2331_o; //(module output)
  assign ctrl_o_rf_rd = n2332_o; //(module output)
  assign ctrl_o_rf_mux = n2333_o; //(module output)
  assign ctrl_o_rf_zero_we = n2334_o; //(module output)
  assign ctrl_o_alu_op = n2335_o; //(module output)
  assign ctrl_o_alu_opa_mux = n2336_o; //(module output)
  assign ctrl_o_alu_opb_mux = n2337_o; //(module output)
  assign ctrl_o_alu_unsigned = n2338_o; //(module output)
  assign ctrl_o_alu_cp_trig = n2339_o; //(module output)
  assign ctrl_o_lsu_req = n2340_o; //(module output)
  assign ctrl_o_lsu_rw = n2341_o; //(module output)
  assign ctrl_o_lsu_mo_we = n2342_o; //(module output)
  assign ctrl_o_lsu_fence = n2343_o; //(module output)
  assign ctrl_o_lsu_priv = n2344_o; //(module output)
  assign ctrl_o_ir_funct3 = n2345_o; //(module output)
  assign ctrl_o_ir_funct12 = n2346_o; //(module output)
  assign ctrl_o_ir_opcode = n2347_o; //(module output)
  assign ctrl_o_cpu_priv = n2348_o; //(module output)
  assign ctrl_o_cpu_sleep = n2349_o; //(module output)
  assign ctrl_o_cpu_trap = n2350_o; //(module output)
  assign ctrl_o_cpu_debug = n2351_o; //(module output)
  assign bus_req_o_addr = n2353_o; //(module output)
  assign bus_req_o_data = n2354_o; //(module output)
  assign bus_req_o_ben = n2355_o; //(module output)
  assign bus_req_o_stb = n2356_o; //(module output)
  assign bus_req_o_rw = n2357_o; //(module output)
  assign bus_req_o_src = n2358_o; //(module output)
  assign bus_req_o_priv = n2359_o; //(module output)
  assign bus_req_o_rvso = n2360_o; //(module output)
  assign bus_req_o_fence = n2361_o; //(module output)
  assign imm_o = n6293_q; //(module output)
  assign fetch_pc_o = n2445_o; //(module output)
  assign curr_pc_o = n2917_o; //(module output)
  assign link_pc_o = n2920_o; //(module output)
  assign csr_rdata_o = n5926_o; //(module output)
  assign xcsr_we_o = n4906_o; //(module output)
  assign xcsr_addr_o = n4907_o; //(module output)
  assign xcsr_wdata_o = n4908_o; //(module output)
  assign n2328_o = n6291_o[0]; // extract
  assign n2329_o = n6291_o[5:1]; // extract
  assign n2330_o = n6291_o[10:6]; // extract
  assign n2331_o = n6291_o[15:11]; // extract
  assign n2332_o = n6291_o[20:16]; // extract
  assign n2333_o = n6291_o[22:21]; // extract
  assign n2334_o = n6291_o[23]; // extract
  assign n2335_o = n6291_o[26:24]; // extract
  assign n2336_o = n6291_o[27]; // extract
  assign n2337_o = n6291_o[28]; // extract
  assign n2338_o = n6291_o[29]; // extract
  assign n2339_o = n6291_o[35:30]; // extract
  assign n2340_o = n6291_o[36]; // extract
  assign n2341_o = n6291_o[37]; // extract
  assign n2342_o = n6291_o[38]; // extract
  assign n2343_o = n6291_o[39]; // extract
  assign n2344_o = n6291_o[40]; // extract
  assign n2345_o = n6291_o[43:41]; // extract
  assign n2346_o = n6291_o[55:44]; // extract
  assign n2347_o = n6291_o[62:56]; // extract
  assign n2348_o = n6291_o[63]; // extract
  assign n2349_o = n6291_o[64]; // extract
  assign n2350_o = n6291_o[65]; // extract
  assign n2351_o = n6291_o[66]; // extract
  assign n2353_o = n6292_o[31:0]; // extract
  assign n2354_o = n6292_o[63:32]; // extract
  assign n2355_o = n6292_o[67:64]; // extract
  assign n2356_o = n6292_o[68]; // extract
  assign n2357_o = n6292_o[69]; // extract
  assign n2358_o = n6292_o[70]; // extract
  assign n2359_o = n6292_o[71]; // extract
  assign n2360_o = n6292_o[72]; // extract
  assign n2361_o = n6292_o[73]; // extract
  assign n2362_o = {bus_rsp_i_err, bus_rsp_i_ack, bus_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:142:10  */
  assign fetch_engine = n6238_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:151:10  */
  assign ipb = n6239_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:164:10  */
  assign issue_engine = n6241_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:180:10  */
  assign decode_aux = n6242_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:200:10  */
  assign execute_engine = n6253_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:208:10  */
  assign monitor = n6255_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:211:10  */
  assign sleep_mode = n6256_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:235:10  */
  assign trap_ctrl = n6261_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:238:10  */
  assign ctrl = n6262_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:238:16  */
  assign ctrl_nxt = n6263_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:290:10  */
  assign csr = n6273_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:312:10  */
  assign cnt = n6285_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:313:10  */
  assign cnt_lo_rd = n6286_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:314:10  */
  assign cnt_hi_rd = n6287_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:317:10  */
  assign cnt_event = n6288_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:327:10  */
  assign debug_ctrl = n6289_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:330:10  */
  assign illegal_cmd = n4185_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:333:10  */
  assign csr_reg_valid = n3858_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:334:10  */
  assign csr_rw_valid = n3877_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:335:10  */
  assign csr_priv_valid = n3914_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:338:28  */
  assign hw_trigger_fired = 1'b0; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:341:10  */
  assign csr_rdata = n6290_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:341:21  */
  assign xcsr_rdata = xcsr_rdata_i; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:353:16  */
  assign n2372_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:360:24  */
  assign n2378_o = fetch_engine[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:360:30  */
  assign n2380_o = n2378_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:363:46  */
  assign n2382_o = fetch_engine[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:363:70  */
  assign n2383_o = fetch_engine[35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:363:54  */
  assign n2384_o = n2382_o | n2383_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:360:7  */
  assign n2385_o = n2380_o ? 1'b0 : n2384_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:367:25  */
  assign n2386_o = fetch_engine[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:371:19  */
  assign n2387_o = ipb[73:72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:371:24  */
  assign n2389_o = n2387_o == 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:373:31  */
  assign n2391_o = fetch_engine[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:373:63  */
  assign n2392_o = fetch_engine[35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:373:46  */
  assign n2393_o = n2391_o | n2392_o;
  assign n2395_o = fetch_engine[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:373:11  */
  assign n2396_o = n2393_o ? 2'b00 : n2395_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:371:11  */
  assign n2397_o = n2389_o ? 2'b10 : n2396_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:369:9  */
  assign n2399_o = n2386_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:379:28  */
  assign n2400_o = fetch_engine[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:380:75  */
  assign n2401_o = fetch_engine[34:3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:380:79  */
  assign n2403_o = n2401_o + 32'b00000000000000000000000000000100;
  assign n2405_o = n2403_o[31:2]; // extract
  assign n2406_o = n2403_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:382:30  */
  assign n2407_o = fetch_engine[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:382:62  */
  assign n2408_o = fetch_engine[35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:382:45  */
  assign n2409_o = n2407_o | n2408_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:382:13  */
  assign n2412_o = n2409_o ? 2'b00 : 2'b01;
  assign n2413_o = {n2405_o, 1'b0, n2406_o};
  assign n2414_o = fetch_engine[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:379:11  */
  assign n2415_o = n2400_o ? n2412_o : n2414_o;
  assign n2416_o = fetch_engine[34:3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:379:11  */
  assign n2417_o = n2400_o ? n2413_o : n2416_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:377:9  */
  assign n2419_o = n2386_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:391:55  */
  assign n2420_o = execute_engine[139:109]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:391:73  */
  assign n2422_o = {n2420_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:392:37  */
  assign n2423_o = csr[153]; // extract
  assign n2425_o = {n2419_o, n2399_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:367:7  */
  always @*
    case (n2425_o)
      2'b10: n2426_o = n2415_o;
      2'b01: n2426_o = n2397_o;
      default: n2426_o = 2'b01;
    endcase
  assign n2427_o = fetch_engine[34:3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:367:7  */
  always @*
    case (n2425_o)
      2'b10: n2428_o = n2417_o;
      2'b01: n2428_o = n2427_o;
      default: n2428_o = n2422_o;
    endcase
  assign n2429_o = fetch_engine[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:367:7  */
  always @*
    case (n2425_o)
      2'b10: n2430_o = n2429_o;
      2'b01: n2430_o = n2429_o;
      default: n2430_o = n2423_o;
    endcase
  assign n2431_o = {n2428_o, n2385_o, n2426_o};
  assign n2436_o = {32'b00000000000000000000000000000000, 1'b1, 2'b00};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:400:36  */
  assign n2440_o = fetch_engine[34:5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:400:54  */
  assign n2442_o = {n2440_o, 2'b00};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:401:36  */
  assign n2443_o = fetch_engine[34:5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:401:54  */
  assign n2445_o = {n2443_o, 2'b00};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:404:43  */
  assign n2447_o = fetch_engine[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:404:49  */
  assign n2449_o = n2447_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:404:72  */
  assign n2450_o = ipb[73:72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:404:77  */
  assign n2452_o = n2450_o == 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:404:63  */
  assign n2453_o = n2452_o & n2449_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:404:24  */
  assign n2454_o = n2453_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:407:34  */
  assign n2456_o = n2362_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:407:51  */
  assign n2457_o = n2362_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:407:38  */
  assign n2458_o = n2456_o | n2457_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:410:30  */
  assign n2459_o = n2362_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:410:34  */
  assign n2460_o = n2459_o | i_pmp_fault_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:410:68  */
  assign n2461_o = n2362_o[15:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:410:52  */
  assign n2462_o = {n2460_o, n2461_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:411:30  */
  assign n2463_o = n2362_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:411:34  */
  assign n2464_o = n2463_o | i_pmp_fault_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:411:68  */
  assign n2465_o = n2362_o[31:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:411:52  */
  assign n2466_o = {n2464_o, n2465_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:414:39  */
  assign n2468_o = fetch_engine[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:414:45  */
  assign n2470_o = n2468_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:414:77  */
  assign n2471_o = fetch_engine[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:414:59  */
  assign n2472_o = n2471_o & n2470_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:415:42  */
  assign n2473_o = fetch_engine[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:415:46  */
  assign n2474_o = ~n2473_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:415:53  */
  assign n2476_o = n2474_o | 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:414:89  */
  assign n2477_o = n2476_o & n2472_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:414:20  */
  assign n2478_o = n2477_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:416:39  */
  assign n2481_o = fetch_engine[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:416:45  */
  assign n2483_o = n2481_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:416:77  */
  assign n2484_o = fetch_engine[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:416:59  */
  assign n2485_o = n2484_o & n2483_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:416:20  */
  assign n2486_o = n2485_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:419:35  */
  assign n2488_o = fetch_engine[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:425:27  */
  assign n2494_o = ctrl[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:432:5  */
  neorv32_fifo_2_17_29e2dcfbb16f63bb0254df7585a15bb6fb5e927d prefetch_buffer_n1_prefetch_buffer_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n2495_o),
    .wdata_i(n2496_o),
    .we_i(n2497_o),
    .re_i(n2499_o),
    .half_o(),
    .free_o(prefetch_buffer_n1_prefetch_buffer_inst_free_o),
    .rdata_o(prefetch_buffer_n1_prefetch_buffer_inst_rdata_o),
    .avail_o(prefetch_buffer_n1_prefetch_buffer_inst_avail_o));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:444:31  */
  assign n2495_o = fetch_engine[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:447:27  */
  assign n2496_o = ipb[33:17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:448:24  */
  assign n2497_o = ipb[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:451:24  */
  assign n2499_o = ipb[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:432:5  */
  neorv32_fifo_2_17_29e2dcfbb16f63bb0254df7585a15bb6fb5e927d prefetch_buffer_n2_prefetch_buffer_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n2502_o),
    .wdata_i(n2503_o),
    .we_i(n2504_o),
    .re_i(n2506_o),
    .half_o(),
    .free_o(prefetch_buffer_n2_prefetch_buffer_inst_free_o),
    .rdata_o(prefetch_buffer_n2_prefetch_buffer_inst_rdata_o),
    .avail_o(prefetch_buffer_n2_prefetch_buffer_inst_avail_o));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:444:31  */
  assign n2502_o = fetch_engine[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:447:27  */
  assign n2503_o = ipb[16:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:448:24  */
  assign n2504_o = ipb[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:451:24  */
  assign n2506_o = ipb[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:466:5  */
  neorv32_cpu_decompressor neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst (
    .ci_instr16_i(n2509_o),
    .ci_instr32_o(neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_instr32_o));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:468:36  */
  assign n2509_o = issue_engine[18:3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:479:38  */
  assign n2511_o = ipb[66:51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:479:71  */
  assign n2512_o = issue_engine[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:479:77  */
  assign n2513_o = ~n2512_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:479:52  */
  assign n2514_o = n2513_o ? n2511_o : n2515_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:479:101  */
  assign n2515_o = ipb[49:34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:489:18  */
  assign n2517_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:492:26  */
  assign n2520_o = fetch_engine[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:493:55  */
  assign n2521_o = execute_engine[109]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:494:29  */
  assign n2522_o = issue_engine[87]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:495:47  */
  assign n2523_o = issue_engine[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:495:75  */
  assign n2524_o = issue_engine[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:495:58  */
  assign n2525_o = ~n2524_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:495:53  */
  assign n2526_o = n2523_o & n2525_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:495:103  */
  assign n2527_o = issue_engine[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:495:87  */
  assign n2528_o = n2526_o | n2527_o;
  assign n2529_o = issue_engine[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:494:9  */
  assign n2530_o = n2522_o ? n2528_o : n2529_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:492:9  */
  assign n2531_o = n2520_o ? n2521_o : n2530_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:507:24  */
  assign n2540_o = issue_engine[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:507:30  */
  assign n2541_o = ~n2540_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:508:25  */
  assign n2542_o = ipb[52:51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:508:38  */
  assign n2544_o = n2542_o != 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:509:46  */
  assign n2545_o = ipb[74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:510:46  */
  assign n2546_o = ipb[74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:511:55  */
  assign n2547_o = ipb[67]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:511:41  */
  assign n2549_o = {1'b1, n2547_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:511:75  */
  assign n2550_o = issue_engine[50:19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:511:60  */
  assign n2551_o = {n2549_o, n2550_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:513:54  */
  assign n2552_o = ipb[74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:513:71  */
  assign n2553_o = ipb[75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:513:58  */
  assign n2554_o = n2552_o & n2553_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:513:54  */
  assign n2555_o = ipb[74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:513:71  */
  assign n2556_o = ipb[75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:513:58  */
  assign n2557_o = n2555_o & n2556_o;
  assign n2558_o = {n2554_o, n2557_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:514:51  */
  assign n2559_o = ipb[67]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:514:37  */
  assign n2561_o = {1'b0, n2559_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:514:70  */
  assign n2562_o = ipb[49:34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:514:56  */
  assign n2563_o = {n2561_o, n2562_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:514:98  */
  assign n2564_o = ipb[66:51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:514:84  */
  assign n2565_o = {n2563_o, n2564_o};
  assign n2566_o = {n2558_o, n2565_o};
  assign n2567_o = {n2546_o, n2551_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:507:7  */
  assign n2568_o = n2609_o ? n2545_o : 1'b0;
  assign n2569_o = n2566_o[34:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:508:9  */
  assign n2570_o = n2544_o ? n2567_o : n2569_o;
  assign n2571_o = n2566_o[35]; // extract
  assign n2572_o = n2539_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:508:9  */
  assign n2573_o = n2544_o ? n2572_o : n2571_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:518:25  */
  assign n2574_o = ipb[35:34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:518:38  */
  assign n2576_o = n2574_o != 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:519:46  */
  assign n2577_o = ipb[75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:520:46  */
  assign n2578_o = ipb[75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:521:55  */
  assign n2579_o = ipb[50]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:521:41  */
  assign n2581_o = {1'b1, n2579_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:521:75  */
  assign n2582_o = issue_engine[50:19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:521:60  */
  assign n2583_o = {n2581_o, n2582_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:523:54  */
  assign n2584_o = ipb[74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:523:71  */
  assign n2585_o = ipb[75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:523:58  */
  assign n2586_o = n2584_o & n2585_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:523:54  */
  assign n2587_o = ipb[74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:523:71  */
  assign n2588_o = ipb[75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:523:58  */
  assign n2589_o = n2587_o & n2588_o;
  assign n2590_o = {n2586_o, n2589_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:524:51  */
  assign n2591_o = ipb[67]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:524:37  */
  assign n2593_o = {1'b0, n2591_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:524:70  */
  assign n2594_o = ipb[66:51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:524:56  */
  assign n2595_o = {n2593_o, n2594_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:524:98  */
  assign n2596_o = ipb[49:34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:524:84  */
  assign n2597_o = {n2595_o, n2596_o};
  assign n2598_o = {n2590_o, n2597_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:518:9  */
  assign n2599_o = n2576_o ? n2577_o : 1'b0;
  assign n2600_o = n2598_o[33:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:518:9  */
  assign n2601_o = n2576_o ? n2583_o : n2600_o;
  assign n2602_o = n2598_o[34]; // extract
  assign n2603_o = n2539_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:518:9  */
  assign n2604_o = n2576_o ? n2603_o : n2602_o;
  assign n2605_o = n2598_o[35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:518:9  */
  assign n2606_o = n2576_o ? n2578_o : n2605_o;
  assign n2607_o = {n2606_o, n2604_o, n2601_o};
  assign n2608_o = {n2573_o, n2570_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:507:7  */
  assign n2609_o = n2544_o & n2541_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:507:7  */
  assign n2610_o = n2541_o ? 1'b0 : n2599_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:507:7  */
  assign n2611_o = n2541_o ? n2608_o : n2607_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:538:34  */
  assign n2613_o = issue_engine[85]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:538:55  */
  assign n2614_o = issue_engine[87]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:538:38  */
  assign n2615_o = n2613_o & n2614_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:539:34  */
  assign n2616_o = issue_engine[86]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:539:55  */
  assign n2617_o = issue_engine[87]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:539:38  */
  assign n2618_o = n2616_o & n2617_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:550:16  */
  assign n2620_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2622_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2623_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2624_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2625_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2626_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2627_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2628_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2629_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2630_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2631_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2632_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2633_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2634_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2635_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2636_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2637_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2638_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2639_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2640_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2641_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:554:62  */
  assign n2642_o = execute_engine[39]; // extract
  assign n2643_o = {n2622_o, n2623_o, n2624_o, n2625_o};
  assign n2644_o = {n2626_o, n2627_o, n2628_o, n2629_o};
  assign n2645_o = {n2630_o, n2631_o, n2632_o, n2633_o};
  assign n2646_o = {n2634_o, n2635_o, n2636_o, n2637_o};
  assign n2647_o = {n2638_o, n2639_o, n2640_o, n2641_o};
  assign n2648_o = {n2643_o, n2644_o, n2645_o, n2646_o};
  assign n2649_o = {n2647_o, n2642_o};
  assign n2650_o = {n2648_o, n2649_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:556:51  */
  assign n2652_o = execute_engine[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:558:23  */
  assign n2653_o = decode_aux[6:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2654_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2655_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2656_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2657_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2658_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2659_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2660_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2661_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2662_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2663_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2664_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2665_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2666_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2667_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2668_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2669_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2670_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2671_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2672_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2673_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:560:66  */
  assign n2674_o = execute_engine[39]; // extract
  assign n2675_o = {n2654_o, n2655_o, n2656_o, n2657_o};
  assign n2676_o = {n2658_o, n2659_o, n2660_o, n2661_o};
  assign n2677_o = {n2662_o, n2663_o, n2664_o, n2665_o};
  assign n2678_o = {n2666_o, n2667_o, n2668_o, n2669_o};
  assign n2679_o = {n2670_o, n2671_o, n2672_o, n2673_o};
  assign n2680_o = {n2675_o, n2676_o, n2677_o, n2678_o};
  assign n2681_o = {n2679_o, n2674_o};
  assign n2682_o = {n2680_o, n2681_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:561:55  */
  assign n2683_o = execute_engine[38:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:562:55  */
  assign n2684_o = execute_engine[19:15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:559:9  */
  assign n2686_o = n2653_o == 7'b0100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2687_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2688_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2689_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2690_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2691_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2692_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2693_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2694_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2695_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2696_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2697_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2698_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2699_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2700_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2701_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2702_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2703_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2704_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2705_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:564:66  */
  assign n2706_o = execute_engine[39]; // extract
  assign n2707_o = {n2687_o, n2688_o, n2689_o, n2690_o};
  assign n2708_o = {n2691_o, n2692_o, n2693_o, n2694_o};
  assign n2709_o = {n2695_o, n2696_o, n2697_o, n2698_o};
  assign n2710_o = {n2699_o, n2700_o, n2701_o, n2702_o};
  assign n2711_o = {n2703_o, n2704_o, n2705_o, n2706_o};
  assign n2712_o = {n2707_o, n2708_o, n2709_o, n2710_o};
  assign n2713_o = {n2712_o, n2711_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:565:55  */
  assign n2714_o = execute_engine[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:566:55  */
  assign n2715_o = execute_engine[38:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:567:55  */
  assign n2716_o = execute_engine[19:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:563:9  */
  assign n2719_o = n2653_o == 7'b1100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:570:55  */
  assign n2720_o = execute_engine[39:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:569:9  */
  assign n2723_o = n2653_o == 7'b0110111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:569:27  */
  assign n2725_o = n2653_o == 7'b0010111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:569:27  */
  assign n2726_o = n2723_o | n2725_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2727_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2728_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2729_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2730_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2731_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2732_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2733_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2734_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2735_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2736_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2737_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:573:66  */
  assign n2738_o = execute_engine[39]; // extract
  assign n2739_o = {n2727_o, n2728_o, n2729_o, n2730_o};
  assign n2740_o = {n2731_o, n2732_o, n2733_o, n2734_o};
  assign n2741_o = {n2735_o, n2736_o, n2737_o, n2738_o};
  assign n2742_o = {n2739_o, n2740_o, n2741_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:574:55  */
  assign n2743_o = execute_engine[27:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:575:55  */
  assign n2744_o = execute_engine[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:576:55  */
  assign n2745_o = execute_engine[38:29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:572:9  */
  assign n2748_o = n2653_o == 7'b1101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:578:9  */
  assign n2750_o = n2653_o == 7'b0101111;
  assign n2751_o = {n2750_o, n2748_o, n2726_o, n2719_o, n2686_o};
  assign n2752_o = n2684_o[0]; // extract
  assign n2753_o = n2721_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:558:7  */
  always @*
    case (n2751_o)
      5'b10000: n2754_o = n2652_o;
      5'b01000: n2754_o = 1'b0;
      5'b00100: n2754_o = n2753_o;
      5'b00010: n2754_o = 1'b0;
      5'b00001: n2754_o = n2752_o;
      default: n2754_o = n2652_o;
    endcase
  assign n2755_o = n2684_o[4:1]; // extract
  assign n2756_o = n2721_o[4:1]; // extract
  assign n2757_o = n2745_o[3:0]; // extract
  assign n2758_o = execute_engine[32:29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:558:7  */
  always @*
    case (n2751_o)
      5'b10000: n2759_o = n2758_o;
      5'b01000: n2759_o = n2757_o;
      5'b00100: n2759_o = n2756_o;
      5'b00010: n2759_o = n2716_o;
      5'b00001: n2759_o = n2755_o;
      default: n2759_o = n2758_o;
    endcase
  assign n2760_o = n2721_o[10:5]; // extract
  assign n2761_o = n2745_o[9:4]; // extract
  assign n2762_o = execute_engine[38:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:558:7  */
  always @*
    case (n2751_o)
      5'b10000: n2763_o = n2762_o;
      5'b01000: n2763_o = n2761_o;
      5'b00100: n2763_o = n2760_o;
      5'b00010: n2763_o = n2715_o;
      5'b00001: n2763_o = n2683_o;
      default: n2763_o = n2762_o;
    endcase
  assign n2764_o = n2682_o[0]; // extract
  assign n2765_o = n2721_o[11]; // extract
  assign n2766_o = n2650_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:558:7  */
  always @*
    case (n2751_o)
      5'b10000: n2767_o = n2766_o;
      5'b01000: n2767_o = n2744_o;
      5'b00100: n2767_o = n2765_o;
      5'b00010: n2767_o = n2714_o;
      5'b00001: n2767_o = n2764_o;
      default: n2767_o = n2766_o;
    endcase
  assign n2768_o = n2682_o[8:1]; // extract
  assign n2769_o = n2713_o[7:0]; // extract
  assign n2770_o = n2720_o[7:0]; // extract
  assign n2771_o = n2650_o[8:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:558:7  */
  always @*
    case (n2751_o)
      5'b10000: n2772_o = n2771_o;
      5'b01000: n2772_o = n2743_o;
      5'b00100: n2772_o = n2770_o;
      5'b00010: n2772_o = n2769_o;
      5'b00001: n2772_o = n2768_o;
      default: n2772_o = n2771_o;
    endcase
  assign n2773_o = n2682_o[20:9]; // extract
  assign n2774_o = n2713_o[19:8]; // extract
  assign n2775_o = n2720_o[19:8]; // extract
  assign n2776_o = n2650_o[20:9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:558:7  */
  always @*
    case (n2751_o)
      5'b10000: n2777_o = n2776_o;
      5'b01000: n2777_o = n2742_o;
      5'b00100: n2777_o = n2775_o;
      5'b00010: n2777_o = n2774_o;
      5'b00001: n2777_o = n2773_o;
      default: n2777_o = n2776_o;
    endcase
  assign n2781_o = {n2777_o, n2772_o, n2767_o, n2763_o, n2759_o, n2754_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:595:26  */
  assign n2787_o = execute_engine[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:595:49  */
  assign n2788_o = ~n2787_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:596:28  */
  assign n2789_o = execute_engine[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:596:49  */
  assign n2790_o = ~n2789_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:597:45  */
  assign n2791_o = cmp_i[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:597:80  */
  assign n2792_o = execute_engine[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:597:59  */
  assign n2793_o = n2791_o ^ n2792_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:599:45  */
  assign n2794_o = cmp_i[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:599:79  */
  assign n2795_o = execute_engine[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:599:58  */
  assign n2796_o = n2794_o ^ n2795_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:596:7  */
  assign n2797_o = n2790_o ? n2793_o : n2796_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:595:5  */
  assign n2799_o = n2788_o ? n2797_o : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:611:16  */
  assign n2802_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:624:46  */
  assign n2810_o = execute_engine[7:4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:625:46  */
  assign n2811_o = execute_engine[71:40]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:626:46  */
  assign n2812_o = execute_engine[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:629:26  */
  assign n2813_o = execute_engine[107]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:630:52  */
  assign n2814_o = execute_engine[139:109]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:630:70  */
  assign n2816_o = {n2814_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:634:26  */
  assign n2819_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:634:32  */
  assign n2821_o = n2819_o == 4'b1000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:635:57  */
  assign n2822_o = execute_engine[139:109]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:635:75  */
  assign n2824_o = {n2822_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:639:27  */
  assign n2827_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:647:26  */
  assign n2830_o = csr[193:192]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:647:39  */
  assign n2832_o = n2830_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:647:67  */
  assign n2833_o = trap_ctrl[61]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:647:47  */
  assign n2834_o = n2833_o & n2832_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:648:50  */
  assign n2835_o = csr[223:199]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:648:85  */
  assign n2836_o = trap_ctrl[59:55]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:648:68  */
  assign n2837_o = {n2835_o, n2836_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:648:98  */
  assign n2839_o = {n2837_o, 2'b00};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:650:50  */
  assign n2840_o = csr[223:194]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:650:68  */
  assign n2842_o = {n2840_o, 2'b00};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:647:13  */
  assign n2843_o = n2834_o ? n2839_o : n2842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:641:9  */
  assign n2845_o = n2827_o == 4'b0001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:658:47  */
  assign n2847_o = csr[185:155]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:658:65  */
  assign n2849_o = {n2847_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:654:9  */
  assign n2851_o = n2827_o == 4'b0010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:662:32  */
  assign n2852_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:662:48  */
  assign n2853_o = ~n2852_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:662:75  */
  assign n2854_o = execute_engine[74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:662:55  */
  assign n2855_o = n2854_o & n2853_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:663:48  */
  assign n2856_o = alu_add_i[31:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:663:66  */
  assign n2858_o = {n2856_o, 1'b0};
  assign n2859_o = execute_engine[139:108]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:662:11  */
  assign n2860_o = n2855_o ? n2858_o : n2859_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:661:9  */
  assign n2862_o = n2827_o == 4'b1000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:667:79  */
  assign n2863_o = execute_engine[106:75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:667:109  */
  assign n2864_o = execute_engine[171:140]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:667:83  */
  assign n2865_o = n2863_o + n2864_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:666:9  */
  assign n2867_o = n2827_o == 4'b0110;
  assign n2868_o = {n2867_o, n2862_o, n2851_o, n2845_o};
  assign n2869_o = execute_engine[139:108]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:639:7  */
  always @*
    case (n2868_o)
      4'b1000: n2870_o = n2865_o;
      4'b0100: n2870_o = n2860_o;
      4'b0010: n2870_o = n2849_o;
      4'b0001: n2870_o = n2843_o;
      default: n2870_o = n2869_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:677:29  */
  assign n2905_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:683:72  */
  assign n2909_o = execute_engine[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:683:78  */
  assign n2910_o = ~n2909_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:683:85  */
  assign n2912_o = n2910_o | 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:683:50  */
  assign n2913_o = n2912_o ? 4'b0100 : 4'b0010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:686:33  */
  assign n2915_o = execute_engine[106:76]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:686:51  */
  assign n2917_o = {n2915_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:687:38  */
  assign n2918_o = execute_engine[203:173]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:687:56  */
  assign n2920_o = {n2918_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:769:26  */
  assign n2930_o = execute_engine[39:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:769:73  */
  assign n2932_o = n2930_o == 7'b0000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:770:103  */
  assign n2933_o = execute_engine[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:770:124  */
  assign n2934_o = ~n2933_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:770:81  */
  assign n2936_o = n2934_o & 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:770:7  */
  assign n2938_o = n2936_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:773:63  */
  assign n2939_o = execute_engine[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:773:41  */
  assign n2941_o = n2939_o & 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:773:7  */
  assign n2943_o = n2941_o ? 1'b1 : 1'b0;
  assign n2944_o = {n2943_o, n2938_o};
  assign n2945_o = {1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:769:5  */
  assign n2946_o = n2932_o ? n2944_o : n2945_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:786:53  */
  assign n2949_o = execute_engine[27:23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:786:94  */
  assign n2951_o = n2949_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:786:30  */
  assign n2952_o = n2951_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:787:53  */
  assign n2955_o = execute_engine[19:15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:787:94  */
  assign n2957_o = n2955_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:787:30  */
  assign n2958_o = n2957_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:790:41  */
  assign n2960_o = execute_engine[14:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:790:90  */
  assign n2962_o = {n2960_o, 2'b11};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:798:48  */
  assign n2964_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:799:48  */
  assign n2965_o = execute_engine[39:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:800:48  */
  assign n2966_o = execute_engine[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:820:26  */
  assign n2978_o = execute_engine[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:821:49  */
  assign n2979_o = execute_engine[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:823:49  */
  assign n2980_o = execute_engine[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:820:5  */
  assign n2981_o = n2978_o ? n2979_o : n2980_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:827:21  */
  assign n2985_o = decode_aux[6:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:828:7  */
  assign n2988_o = n2985_o == 7'b0010111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:828:27  */
  assign n2990_o = n2985_o == 7'b1101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:828:27  */
  assign n2991_o = n2988_o | n2990_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:828:42  */
  assign n2993_o = n2985_o == 7'b1100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:828:42  */
  assign n2994_o = n2991_o | n2993_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:827:5  */
  always @*
    case (n2994_o)
      1'b1: n2996_o = 1'b1;
      default: n2996_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:835:21  */
  assign n2999_o = decode_aux[6:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:7  */
  assign n3002_o = n2999_o == 7'b0010011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:26  */
  assign n3004_o = n2999_o == 7'b0110111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:26  */
  assign n3005_o = n3002_o | n3004_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:41  */
  assign n3007_o = n2999_o == 7'b0010111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:41  */
  assign n3008_o = n3005_o | n3007_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:58  */
  assign n3010_o = n2999_o == 7'b0000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:58  */
  assign n3011_o = n3008_o | n3010_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:74  */
  assign n3013_o = n2999_o == 7'b0100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:74  */
  assign n3014_o = n3011_o | n3013_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:91  */
  assign n3016_o = n2999_o == 7'b0101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:91  */
  assign n3017_o = n3014_o | n3016_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:106  */
  assign n3019_o = n2999_o == 7'b1100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:106  */
  assign n3020_o = n3017_o | n3019_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:124  */
  assign n3022_o = n2999_o == 7'b1101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:124  */
  assign n3023_o = n3020_o | n3022_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:139  */
  assign n3025_o = n2999_o == 7'b1100111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:836:139  */
  assign n3026_o = n3023_o | n3025_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:835:5  */
  always @*
    case (n3026_o)
      1'b1: n3028_o = 1'b1;
      default: n3028_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:846:43  */
  assign n3029_o = execute_engine[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:25  */
  assign n3032_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:23  */
  assign n3033_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:56  */
  assign n3034_o = trap_ctrl[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:42  */
  assign n3035_o = n3033_o | n3034_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:34  */
  assign n3037_o = issue_engine[85]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:67  */
  assign n3038_o = issue_engine[86]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:45  */
  assign n3039_o = n3037_o | n3038_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:862:56  */
  assign n3041_o = issue_engine[83]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:863:56  */
  assign n3042_o = issue_engine[84]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:864:56  */
  assign n3043_o = issue_engine[82:51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:9  */
  assign n3046_o = n3039_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:9  */
  assign n3047_o = n3039_o ? 4'b0110 : n2964_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:9  */
  assign n3048_o = n3039_o ? n3043_o : n2965_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:9  */
  assign n3049_o = n3039_o ? n3042_o : n2966_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:9  */
  assign n3050_o = n3039_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:860:9  */
  assign n3051_o = n3039_o ? n3041_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:9  */
  assign n3052_o = n3035_o ? 1'b0 : n3046_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:9  */
  assign n3053_o = n3035_o ? 4'b0001 : n3047_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:9  */
  assign n3054_o = n3035_o ? n2965_o : n3048_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:9  */
  assign n3055_o = n3035_o ? n2966_o : n3049_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:9  */
  assign n3056_o = n3035_o ? 1'b0 : n3050_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:854:9  */
  assign n3057_o = n3035_o ? 1'b0 : n3051_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:852:7  */
  assign n3059_o = n3032_o == 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:871:23  */
  assign n3060_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:871:9  */
  assign n3063_o = n3060_o ? 4'b0011 : n2964_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:871:9  */
  assign n3064_o = n3060_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:869:7  */
  assign n3066_o = n3032_o == 4'b0001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:876:7  */
  assign n3070_o = n3032_o == 4'b0010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:881:7  */
  assign n3074_o = n3032_o == 4'b0011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:25  */
  assign n3075_o = decode_aux[6:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:894:35  */
  assign n3076_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:896:39  */
  assign n3077_o = execute_engine[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:896:91  */
  assign n3078_o = execute_engine[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:896:69  */
  assign n3079_o = n3078_o & n3077_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:896:17  */
  assign n3082_o = n3079_o ? 3'b001 : 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:895:15  */
  assign n3084_o = n3076_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:901:15  */
  assign n3087_o = n3076_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:901:33  */
  assign n3089_o = n3076_o == 3'b011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:901:33  */
  assign n3090_o = n3087_o | n3089_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:903:15  */
  assign n3093_o = n3076_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:905:15  */
  assign n3096_o = n3076_o == 3'b110;
  assign n3098_o = {n3096_o, n3093_o, n3090_o, n3084_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:894:13  */
  always @*
    case (n3098_o)
      4'b1000: n3099_o = 3'b110;
      4'b0100: n3099_o = 3'b101;
      4'b0010: n3099_o = 3'b011;
      4'b0001: n3099_o = n3082_o;
      default: n3099_o = 3'b111;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:912:70  */
  assign n3100_o = execute_engine[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:912:48  */
  assign n3102_o = n3100_o & 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:913:30  */
  assign n3103_o = decode_aux[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:913:61  */
  assign n3104_o = decode_aux[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:913:46  */
  assign n3105_o = n3103_o | n3104_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:912:112  */
  assign n3106_o = n3105_o & n3102_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:913:79  */
  assign n3108_o = n3106_o | 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:930:37  */
  assign n3111_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:930:84  */
  assign n3113_o = n3111_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:931:37  */
  assign n3114_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:931:84  */
  assign n3116_o = n3114_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:930:100  */
  assign n3117_o = n3113_o | n3116_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:930:13  */
  assign n3122_o = n3117_o ? 4'b0111 : 4'b0000;
  assign n3123_o = n2982_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:930:13  */
  assign n3124_o = n3117_o ? n3123_o : 1'b1;
  assign n3125_o = n2982_o[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:930:13  */
  assign n3126_o = n3117_o ? 1'b1 : n3125_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:912:13  */
  assign n3127_o = n3108_o ? 4'b0111 : n3122_o;
  assign n3128_o = n2982_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:912:13  */
  assign n3129_o = n3108_o ? n3128_o : n3124_o;
  assign n3130_o = n2982_o[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:912:13  */
  assign n3131_o = n3108_o ? n3130_o : n3126_o;
  assign n3132_o = n2982_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:912:13  */
  assign n3133_o = n3108_o ? 1'b1 : n3132_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:892:11  */
  assign n3135_o = n3075_o == 7'b0110011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:892:29  */
  assign n3137_o = n3075_o == 7'b0010011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:892:29  */
  assign n3138_o = n3135_o | n3137_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:942:34  */
  assign n3139_o = execute_engine[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:942:13  */
  assign n3141_o = n3139_o ? 3'b100 : 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:941:11  */
  assign n3145_o = n3075_o == 7'b0110111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:941:29  */
  assign n3147_o = n3075_o == 7'b0010111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:941:29  */
  assign n3148_o = n3145_o | n3147_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:951:11  */
  assign n3151_o = n3075_o == 7'b0000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:951:30  */
  assign n3153_o = n3075_o == 7'b0100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:951:30  */
  assign n3154_o = n3151_o | n3153_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:951:47  */
  assign n3156_o = n3075_o == 7'b0101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:951:47  */
  assign n3157_o = n3154_o | n3156_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:955:11  */
  assign n3160_o = n3075_o == 7'b1100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:955:32  */
  assign n3162_o = n3075_o == 7'b1101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:955:32  */
  assign n3163_o = n3160_o | n3162_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:955:47  */
  assign n3165_o = n3075_o == 7'b1100111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:955:47  */
  assign n3166_o = n3163_o | n3165_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:959:11  */
  assign n3169_o = n3075_o == 7'b0001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:963:11  */
  assign n3173_o = n3075_o == 7'b1010011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:968:11  */
  assign n3177_o = n3075_o == 7'b0001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:968:31  */
  assign n3179_o = n3075_o == 7'b0101011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:968:31  */
  assign n3180_o = n3177_o | n3179_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:968:48  */
  assign n3182_o = n3075_o == 7'b1011011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:968:48  */
  assign n3183_o = n3180_o | n3182_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:968:65  */
  assign n3185_o = n3075_o == 7'b1111011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:968:65  */
  assign n3186_o = n3183_o | n3185_o;
  assign n3189_o = {n3186_o, n3173_o, n3169_o, n3166_o, n3157_o, n3148_o, n3138_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:9  */
  always @*
    case (n3189_o)
      7'b1000000: n3190_o = 4'b0111;
      7'b0100000: n3190_o = 4'b0111;
      7'b0010000: n3190_o = 4'b0100;
      7'b0001000: n3190_o = 4'b1000;
      7'b0000100: n3190_o = 4'b1011;
      7'b0000010: n3190_o = 4'b0000;
      7'b0000001: n3190_o = n3127_o;
      default: n3190_o = 4'b1010;
    endcase
  assign n3191_o = n2982_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:9  */
  always @*
    case (n3189_o)
      7'b1000000: n3192_o = n3191_o;
      7'b0100000: n3192_o = n3191_o;
      7'b0010000: n3192_o = n3191_o;
      7'b0001000: n3192_o = n3191_o;
      7'b0000100: n3192_o = n3191_o;
      7'b0000010: n3192_o = 1'b1;
      7'b0000001: n3192_o = n3129_o;
      default: n3192_o = n3191_o;
    endcase
  assign n3193_o = n2982_o[26:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:9  */
  always @*
    case (n3189_o)
      7'b1000000: n3194_o = n3193_o;
      7'b0100000: n3194_o = n3193_o;
      7'b0010000: n3194_o = n3193_o;
      7'b0001000: n3194_o = n3193_o;
      7'b0000100: n3194_o = n3193_o;
      7'b0000010: n3194_o = n3141_o;
      7'b0000001: n3194_o = n3099_o;
      default: n3194_o = n3193_o;
    endcase
  assign n3195_o = n2982_o[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:9  */
  always @*
    case (n3189_o)
      7'b1000000: n3196_o = n3195_o;
      7'b0100000: n3196_o = n3195_o;
      7'b0010000: n3196_o = n3195_o;
      7'b0001000: n3196_o = n3195_o;
      7'b0000100: n3196_o = n3195_o;
      7'b0000010: n3196_o = n3195_o;
      7'b0000001: n3196_o = n3131_o;
      default: n3196_o = n3195_o;
    endcase
  assign n3197_o = n2982_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:9  */
  always @*
    case (n3189_o)
      7'b1000000: n3198_o = n3197_o;
      7'b0100000: n3198_o = n3197_o;
      7'b0010000: n3198_o = n3197_o;
      7'b0001000: n3198_o = n3197_o;
      7'b0000100: n3198_o = n3197_o;
      7'b0000010: n3198_o = n3197_o;
      7'b0000001: n3198_o = n3133_o;
      default: n3198_o = n3197_o;
    endcase
  assign n3199_o = n2982_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:9  */
  always @*
    case (n3189_o)
      7'b1000000: n3200_o = n3199_o;
      7'b0100000: n3200_o = 1'b1;
      7'b0010000: n3200_o = n3199_o;
      7'b0001000: n3200_o = n3199_o;
      7'b0000100: n3200_o = n3199_o;
      7'b0000010: n3200_o = n3199_o;
      7'b0000001: n3200_o = n3199_o;
      default: n3200_o = n3199_o;
    endcase
  assign n3201_o = n2982_o[34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:9  */
  always @*
    case (n3189_o)
      7'b1000000: n3202_o = 1'b1;
      7'b0100000: n3202_o = n3201_o;
      7'b0010000: n3202_o = n3201_o;
      7'b0001000: n3202_o = n3201_o;
      7'b0000100: n3202_o = n3201_o;
      7'b0000010: n3202_o = n3201_o;
      7'b0000001: n3202_o = n3201_o;
      default: n3202_o = n3201_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:889:9  */
  always @*
    case (n3189_o)
      7'b1000000: n3203_o = 1'b0;
      7'b0100000: n3203_o = 1'b0;
      7'b0010000: n3203_o = 1'b0;
      7'b0001000: n3203_o = 1'b0;
      7'b0000100: n3203_o = 1'b0;
      7'b0000010: n3203_o = 1'b0;
      7'b0000001: n3203_o = 1'b0;
      default: n3203_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:886:7  */
  assign n3205_o = n3032_o == 4'b0110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:982:55  */
  assign n3207_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:982:34  */
  assign n3208_o = alu_cp_done_i | n3207_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:982:9  */
  assign n3211_o = n3208_o ? 4'b0000 : n2964_o;
  assign n3212_o = n2982_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:982:9  */
  assign n3213_o = n3208_o ? 1'b1 : n3212_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:979:7  */
  assign n3215_o = n3032_o == 4'b0111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:989:30  */
  assign n3216_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:989:9  */
  assign n3220_o = n3216_o ? 4'b0000 : 4'b0011;
  assign n3221_o = n2982_o[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:989:9  */
  assign n3222_o = n3216_o ? n3221_o : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:987:7  */
  assign n3224_o = n3032_o == 4'b0100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:999:47  */
  assign n3226_o = execute_engine[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1000:30  */
  assign n3227_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1000:46  */
  assign n3228_o = ~n3227_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1000:73  */
  assign n3229_o = execute_engine[74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1000:53  */
  assign n3230_o = n3229_o & n3228_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1000:9  */
  assign n3234_o = n3230_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1000:9  */
  assign n3235_o = n3230_o ? 4'b1001 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:996:7  */
  assign n3237_o = n3032_o == 4'b1000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1007:7  */
  assign n3242_o = n3032_o == 4'b1001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1018:30  */
  assign n3243_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1018:9  */
  assign n3247_o = n3243_o ? 4'b0000 : 4'b1100;
  assign n3248_o = n2982_o[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1018:9  */
  assign n3249_o = n3243_o ? n3248_o : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1016:7  */
  assign n3251_o = n3032_o == 4'b1011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1028:24  */
  assign n3253_o = ~lsu_wait_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1029:30  */
  assign n3254_o = trap_ctrl[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1028:31  */
  assign n3255_o = n3253_o | n3254_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1029:74  */
  assign n3256_o = trap_ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1029:53  */
  assign n3257_o = n3255_o | n3256_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1030:30  */
  assign n3258_o = trap_ctrl[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1029:97  */
  assign n3259_o = n3257_o | n3258_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1030:74  */
  assign n3260_o = trap_ctrl[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1030:53  */
  assign n3261_o = n3259_o | n3260_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1032:32  */
  assign n3262_o = execute_engine[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1032:55  */
  assign n3263_o = ~n3262_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1031:92  */
  assign n3265_o = 1'b0 | n3263_o;
  assign n3267_o = n2982_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1028:9  */
  assign n3268_o = n3272_o ? 1'b1 : n3267_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1028:9  */
  assign n3270_o = n3261_o ? 4'b0000 : n2964_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1028:9  */
  assign n3272_o = n3265_o & n3261_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1025:7  */
  assign n3274_o = n3032_o == 4'b1100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1040:23  */
  assign n3275_o = trap_ctrl[97]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1040:9  */
  assign n3277_o = n3275_o ? 4'b0000 : n2964_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1038:7  */
  assign n3279_o = n3032_o == 4'b0101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1048:30  */
  assign n3281_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1048:77  */
  assign n3283_o = n3281_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1049:30  */
  assign n3284_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1049:46  */
  assign n3285_o = ~n3284_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1048:93  */
  assign n3286_o = n3285_o & n3283_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1050:33  */
  assign n3287_o = execute_engine[39:28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1051:13  */
  assign n3290_o = n3287_o == 12'b000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1052:13  */
  assign n3293_o = n3287_o == 12'b000000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1053:13  */
  assign n3296_o = n3287_o == 12'b001100000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1053:33  */
  assign n3298_o = n3287_o == 12'b011110110010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1053:33  */
  assign n3299_o = n3296_o | n3298_o;
  assign n3301_o = {n3299_o, n3293_o, n3290_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1050:11  */
  always @*
    case (n3301_o)
      3'b100: n3302_o = 4'b0010;
      3'b010: n3302_o = 4'b0000;
      3'b001: n3302_o = 4'b0000;
      default: n3302_o = 4'b0101;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1050:11  */
  always @*
    case (n3301_o)
      3'b100: n3303_o = 1'b0;
      3'b010: n3303_o = 1'b0;
      3'b001: n3303_o = 1'b1;
      default: n3303_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1050:11  */
  always @*
    case (n3301_o)
      3'b100: n3304_o = 1'b0;
      3'b010: n3304_o = 1'b1;
      3'b001: n3304_o = 1'b0;
      default: n3304_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1057:32  */
  assign n3305_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1057:79  */
  assign n3307_o = n3305_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1058:32  */
  assign n3308_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1058:79  */
  assign n3310_o = n3308_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1057:97  */
  assign n3311_o = n3307_o | n3310_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1059:26  */
  assign n3312_o = decode_aux[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1059:35  */
  assign n3313_o = ~n3312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1058:98  */
  assign n3314_o = n3311_o | n3313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1057:11  */
  assign n3316_o = n3314_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1048:9  */
  assign n3318_o = n3286_o ? n3302_o : 4'b0000;
  assign n3319_o = {n3304_o, n3303_o};
  assign n3320_o = {1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1048:9  */
  assign n3321_o = n3286_o ? n3319_o : n3320_o;
  assign n3322_o = n2982_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1048:9  */
  assign n3323_o = n3286_o ? n3322_o : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1048:9  */
  assign n3324_o = n3286_o ? 1'b0 : n3316_o;
  assign n3325_o = {n3279_o, n3274_o, n3251_o, n3242_o, n3237_o, n3224_o, n3215_o, n3205_o, n3074_o, n3070_o, n3066_o, n3059_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3326_o = 1'b0;
      12'b010000000000: n3326_o = 1'b0;
      12'b001000000000: n3326_o = 1'b0;
      12'b000100000000: n3326_o = 1'b0;
      12'b000010000000: n3326_o = n3234_o;
      12'b000001000000: n3326_o = 1'b0;
      12'b000000100000: n3326_o = 1'b0;
      12'b000000010000: n3326_o = 1'b0;
      12'b000000001000: n3326_o = 1'b1;
      12'b000000000100: n3326_o = 1'b0;
      12'b000000000010: n3326_o = 1'b0;
      12'b000000000001: n3326_o = 1'b0;
      default: n3326_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3327_o = 1'b0;
      12'b010000000000: n3327_o = 1'b0;
      12'b001000000000: n3327_o = 1'b0;
      12'b000100000000: n3327_o = 1'b0;
      12'b000010000000: n3327_o = 1'b0;
      12'b000001000000: n3327_o = 1'b0;
      12'b000000100000: n3327_o = 1'b0;
      12'b000000010000: n3327_o = 1'b0;
      12'b000000001000: n3327_o = 1'b0;
      12'b000000000100: n3327_o = 1'b0;
      12'b000000000010: n3327_o = 1'b0;
      12'b000000000001: n3327_o = n3052_o;
      default: n3327_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3328_o = n3277_o;
      12'b010000000000: n3328_o = n3270_o;
      12'b001000000000: n3328_o = n3247_o;
      12'b000100000000: n3328_o = 4'b0000;
      12'b000010000000: n3328_o = n3235_o;
      12'b000001000000: n3328_o = n3220_o;
      12'b000000100000: n3328_o = n3211_o;
      12'b000000010000: n3328_o = n3190_o;
      12'b000000001000: n3328_o = 4'b1001;
      12'b000000000100: n3328_o = 4'b0011;
      12'b000000000010: n3328_o = n3063_o;
      12'b000000000001: n3328_o = n3053_o;
      default: n3328_o = n3318_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3329_o = n2965_o;
      12'b010000000000: n3329_o = n2965_o;
      12'b001000000000: n3329_o = n2965_o;
      12'b000100000000: n3329_o = n2965_o;
      12'b000010000000: n3329_o = n2965_o;
      12'b000001000000: n3329_o = n2965_o;
      12'b000000100000: n3329_o = n2965_o;
      12'b000000010000: n3329_o = n2965_o;
      12'b000000001000: n3329_o = n2965_o;
      12'b000000000100: n3329_o = n2965_o;
      12'b000000000010: n3329_o = n2965_o;
      12'b000000000001: n3329_o = n3054_o;
      default: n3329_o = n2965_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3330_o = n2966_o;
      12'b010000000000: n3330_o = n2966_o;
      12'b001000000000: n3330_o = n2966_o;
      12'b000100000000: n3330_o = n2966_o;
      12'b000010000000: n3330_o = n2966_o;
      12'b000001000000: n3330_o = n2966_o;
      12'b000000100000: n3330_o = n2966_o;
      12'b000000010000: n3330_o = n2966_o;
      12'b000000001000: n3330_o = n2966_o;
      12'b000000000100: n3330_o = n2966_o;
      12'b000000000010: n3330_o = n2966_o;
      12'b000000000001: n3330_o = n3055_o;
      default: n3330_o = n2966_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3331_o = 1'b0;
      12'b010000000000: n3331_o = 1'b0;
      12'b001000000000: n3331_o = 1'b0;
      12'b000100000000: n3331_o = 1'b0;
      12'b000010000000: n3331_o = 1'b0;
      12'b000001000000: n3331_o = 1'b0;
      12'b000000100000: n3331_o = 1'b0;
      12'b000000010000: n3331_o = 1'b0;
      12'b000000001000: n3331_o = 1'b0;
      12'b000000000100: n3331_o = 1'b0;
      12'b000000000010: n3331_o = 1'b0;
      12'b000000000001: n3331_o = n3056_o;
      default: n3331_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3332_o = 1'b0;
      12'b010000000000: n3332_o = 1'b0;
      12'b001000000000: n3332_o = 1'b0;
      12'b000100000000: n3332_o = 1'b0;
      12'b000010000000: n3332_o = 1'b0;
      12'b000001000000: n3332_o = 1'b0;
      12'b000000100000: n3332_o = 1'b0;
      12'b000000010000: n3332_o = 1'b0;
      12'b000000001000: n3332_o = 1'b0;
      12'b000000000100: n3332_o = 1'b0;
      12'b000000000010: n3332_o = n3064_o;
      12'b000000000001: n3332_o = 1'b0;
      default: n3332_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3333_o = 1'b0;
      12'b010000000000: n3333_o = 1'b0;
      12'b001000000000: n3333_o = 1'b0;
      12'b000100000000: n3333_o = 1'b0;
      12'b000010000000: n3333_o = 1'b0;
      12'b000001000000: n3333_o = 1'b0;
      12'b000000100000: n3333_o = 1'b0;
      12'b000000010000: n3333_o = 1'b0;
      12'b000000001000: n3333_o = 1'b0;
      12'b000000000100: n3333_o = 1'b1;
      12'b000000000010: n3333_o = 1'b0;
      12'b000000000001: n3333_o = 1'b0;
      default: n3333_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3334_o = 1'b0;
      12'b010000000000: n3334_o = 1'b0;
      12'b001000000000: n3334_o = 1'b0;
      12'b000100000000: n3334_o = 1'b0;
      12'b000010000000: n3334_o = 1'b0;
      12'b000001000000: n3334_o = 1'b0;
      12'b000000100000: n3334_o = 1'b0;
      12'b000000010000: n3334_o = 1'b0;
      12'b000000001000: n3334_o = 1'b0;
      12'b000000000100: n3334_o = 1'b0;
      12'b000000000010: n3334_o = 1'b0;
      12'b000000000001: n3334_o = n3057_o;
      default: n3334_o = 1'b0;
    endcase
  assign n3335_o = {1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3336_o = n3335_o;
      12'b010000000000: n3336_o = n3335_o;
      12'b001000000000: n3336_o = n3335_o;
      12'b000100000000: n3336_o = n3335_o;
      12'b000010000000: n3336_o = n3335_o;
      12'b000001000000: n3336_o = n3335_o;
      12'b000000100000: n3336_o = n3335_o;
      12'b000000010000: n3336_o = n3335_o;
      12'b000000001000: n3336_o = n3335_o;
      12'b000000000100: n3336_o = n3335_o;
      12'b000000000010: n3336_o = n3335_o;
      12'b000000000001: n3336_o = n3335_o;
      default: n3336_o = n3321_o;
    endcase
  assign n3337_o = n2982_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3338_o = n3337_o;
      12'b010000000000: n3338_o = n3268_o;
      12'b001000000000: n3338_o = n3337_o;
      12'b000100000000: n3338_o = n3337_o;
      12'b000010000000: n3338_o = n3226_o;
      12'b000001000000: n3338_o = n3337_o;
      12'b000000100000: n3338_o = n3213_o;
      12'b000000010000: n3338_o = n3192_o;
      12'b000000001000: n3338_o = n3337_o;
      12'b000000000100: n3338_o = n3337_o;
      12'b000000000010: n3338_o = n3337_o;
      12'b000000000001: n3338_o = n3337_o;
      default: n3338_o = n3323_o;
    endcase
  assign n3339_o = n2982_o[22:21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3340_o = n3339_o;
      12'b010000000000: n3340_o = 2'b01;
      12'b001000000000: n3340_o = n3339_o;
      12'b000100000000: n3340_o = 2'b10;
      12'b000010000000: n3340_o = 2'b11;
      12'b000001000000: n3340_o = n3339_o;
      12'b000000100000: n3340_o = n3339_o;
      12'b000000010000: n3340_o = n3339_o;
      12'b000000001000: n3340_o = n3339_o;
      12'b000000000100: n3340_o = n3339_o;
      12'b000000000010: n3340_o = n3339_o;
      12'b000000000001: n3340_o = n3339_o;
      default: n3340_o = 2'b10;
    endcase
  assign n3341_o = n2982_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3342_o = n3341_o;
      12'b010000000000: n3342_o = n3341_o;
      12'b001000000000: n3342_o = n3341_o;
      12'b000100000000: n3342_o = 1'b1;
      12'b000010000000: n3342_o = n3341_o;
      12'b000001000000: n3342_o = n3341_o;
      12'b000000100000: n3342_o = n3341_o;
      12'b000000010000: n3342_o = n3341_o;
      12'b000000001000: n3342_o = n3341_o;
      12'b000000000100: n3342_o = n3341_o;
      12'b000000000010: n3342_o = n3341_o;
      12'b000000000001: n3342_o = n3341_o;
      default: n3342_o = n3341_o;
    endcase
  assign n3343_o = n2982_o[26:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3344_o = n3343_o;
      12'b010000000000: n3344_o = n3343_o;
      12'b001000000000: n3344_o = n3343_o;
      12'b000100000000: n3344_o = n3343_o;
      12'b000010000000: n3344_o = n3343_o;
      12'b000001000000: n3344_o = n3343_o;
      12'b000000100000: n3344_o = 3'b010;
      12'b000000010000: n3344_o = n3194_o;
      12'b000000001000: n3344_o = n3343_o;
      12'b000000000100: n3344_o = n3343_o;
      12'b000000000010: n3344_o = n3343_o;
      12'b000000000001: n3344_o = n3343_o;
      default: n3344_o = n3343_o;
    endcase
  assign n3345_o = n2982_o[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3346_o = n3345_o;
      12'b010000000000: n3346_o = n3345_o;
      12'b001000000000: n3346_o = n3345_o;
      12'b000100000000: n3346_o = n3345_o;
      12'b000010000000: n3346_o = n3345_o;
      12'b000001000000: n3346_o = n3345_o;
      12'b000000100000: n3346_o = n3345_o;
      12'b000000010000: n3346_o = n3196_o;
      12'b000000001000: n3346_o = n3345_o;
      12'b000000000100: n3346_o = n3345_o;
      12'b000000000010: n3346_o = n3345_o;
      12'b000000000001: n3346_o = n3345_o;
      default: n3346_o = n3345_o;
    endcase
  assign n3347_o = n2982_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3348_o = n3347_o;
      12'b010000000000: n3348_o = n3347_o;
      12'b001000000000: n3348_o = n3347_o;
      12'b000100000000: n3348_o = n3347_o;
      12'b000010000000: n3348_o = n3347_o;
      12'b000001000000: n3348_o = n3347_o;
      12'b000000100000: n3348_o = n3347_o;
      12'b000000010000: n3348_o = n3198_o;
      12'b000000001000: n3348_o = n3347_o;
      12'b000000000100: n3348_o = n3347_o;
      12'b000000000010: n3348_o = n3347_o;
      12'b000000000001: n3348_o = n3347_o;
      default: n3348_o = n3347_o;
    endcase
  assign n3349_o = n2982_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3350_o = n3349_o;
      12'b010000000000: n3350_o = n3349_o;
      12'b001000000000: n3350_o = n3349_o;
      12'b000100000000: n3350_o = n3349_o;
      12'b000010000000: n3350_o = n3349_o;
      12'b000001000000: n3350_o = n3349_o;
      12'b000000100000: n3350_o = n3349_o;
      12'b000000010000: n3350_o = n3200_o;
      12'b000000001000: n3350_o = n3349_o;
      12'b000000000100: n3350_o = n3349_o;
      12'b000000000010: n3350_o = n3349_o;
      12'b000000000001: n3350_o = n3349_o;
      default: n3350_o = n3349_o;
    endcase
  assign n3351_o = n2982_o[34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3352_o = n3351_o;
      12'b010000000000: n3352_o = n3351_o;
      12'b001000000000: n3352_o = n3351_o;
      12'b000100000000: n3352_o = n3351_o;
      12'b000010000000: n3352_o = n3351_o;
      12'b000001000000: n3352_o = n3351_o;
      12'b000000100000: n3352_o = n3351_o;
      12'b000000010000: n3352_o = n3202_o;
      12'b000000001000: n3352_o = n3351_o;
      12'b000000000100: n3352_o = n3351_o;
      12'b000000000010: n3352_o = n3351_o;
      12'b000000000001: n3352_o = n3351_o;
      default: n3352_o = n3351_o;
    endcase
  assign n3353_o = n2982_o[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3354_o = n3353_o;
      12'b010000000000: n3354_o = n3353_o;
      12'b001000000000: n3354_o = n3249_o;
      12'b000100000000: n3354_o = n3353_o;
      12'b000010000000: n3354_o = n3353_o;
      12'b000001000000: n3354_o = n3353_o;
      12'b000000100000: n3354_o = n3353_o;
      12'b000000010000: n3354_o = n3353_o;
      12'b000000001000: n3354_o = n3353_o;
      12'b000000000100: n3354_o = n3353_o;
      12'b000000000010: n3354_o = n3353_o;
      12'b000000000001: n3354_o = n3353_o;
      default: n3354_o = n3353_o;
    endcase
  assign n3355_o = n2982_o[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3356_o = n3355_o;
      12'b010000000000: n3356_o = n3355_o;
      12'b001000000000: n3356_o = n3355_o;
      12'b000100000000: n3356_o = n3355_o;
      12'b000010000000: n3356_o = n3355_o;
      12'b000001000000: n3356_o = n3222_o;
      12'b000000100000: n3356_o = n3355_o;
      12'b000000010000: n3356_o = n3355_o;
      12'b000000001000: n3356_o = n3355_o;
      12'b000000000100: n3356_o = n3355_o;
      12'b000000000010: n3356_o = n3355_o;
      12'b000000000001: n3356_o = n3355_o;
      default: n3356_o = n3355_o;
    endcase
  assign n3359_o = n2982_o[20:1]; // extract
  assign n3364_o = n2982_o[32]; // extract
  assign n3366_o = n2982_o[35]; // extract
  assign n3367_o = n2982_o[66:40]; // extract
  assign n3368_o = n2982_o[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3369_o = 1'b0;
      12'b010000000000: n3369_o = 1'b0;
      12'b001000000000: n3369_o = 1'b0;
      12'b000100000000: n3369_o = 1'b0;
      12'b000010000000: n3369_o = 1'b0;
      12'b000001000000: n3369_o = 1'b0;
      12'b000000100000: n3369_o = 1'b0;
      12'b000000010000: n3369_o = 1'b0;
      12'b000000001000: n3369_o = 1'b0;
      12'b000000000100: n3369_o = 1'b0;
      12'b000000000010: n3369_o = 1'b0;
      12'b000000000001: n3369_o = 1'b0;
      default: n3369_o = n3324_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:850:5  */
  always @*
    case (n3325_o)
      12'b100000000000: n3370_o = 1'b0;
      12'b010000000000: n3370_o = 1'b0;
      12'b001000000000: n3370_o = 1'b0;
      12'b000100000000: n3370_o = 1'b0;
      12'b000010000000: n3370_o = 1'b0;
      12'b000001000000: n3370_o = 1'b0;
      12'b000000100000: n3370_o = 1'b0;
      12'b000000010000: n3370_o = n3203_o;
      12'b000000001000: n3370_o = 1'b0;
      12'b000000000100: n3370_o = 1'b0;
      12'b000000000010: n3370_o = 1'b0;
      12'b000000000001: n3370_o = 1'b0;
      default: n3370_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1073:16  */
  assign n3373_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1076:26  */
  assign n3375_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1076:32  */
  assign n3377_o = n3375_o == 4'b0101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1077:15  */
  assign n3378_o = ipb[73:72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1077:20  */
  assign n3380_o = n3378_o != 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1076:41  */
  assign n3381_o = n3380_o & n3377_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1078:21  */
  assign n3382_o = trap_ctrl[97]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1078:28  */
  assign n3383_o = ~n3382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1077:29  */
  assign n3384_o = n3383_o & n3381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1076:7  */
  assign n3387_o = n3384_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1091:31  */
  assign n3392_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1092:48  */
  assign n3393_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1092:27  */
  assign n3394_o = ~n3393_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1091:40  */
  assign n3395_o = n3392_o & n3394_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:48  */
  assign n3396_o = trap_ctrl[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:27  */
  assign n3397_o = ~n3396_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1092:65  */
  assign n3398_o = n3395_o & n3397_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:91  */
  assign n3399_o = trap_ctrl[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:70  */
  assign n3400_o = ~n3399_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:65  */
  assign n3401_o = n3398_o & n3400_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:134  */
  assign n3402_o = trap_ctrl[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:113  */
  assign n3403_o = ~n3402_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:108  */
  assign n3404_o = n3401_o & n3403_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1094:48  */
  assign n3405_o = trap_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1094:27  */
  assign n3406_o = ~n3405_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1093:150  */
  assign n3407_o = n3404_o & n3406_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1094:91  */
  assign n3408_o = trap_ctrl[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1094:70  */
  assign n3409_o = ~n3408_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1094:65  */
  assign n3410_o = n3407_o & n3409_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1094:134  */
  assign n3411_o = trap_ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1094:113  */
  assign n3412_o = ~n3411_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1094:108  */
  assign n3413_o = n3410_o & n3412_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1095:43  */
  assign n3414_o = execute_engine[27:23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1096:43  */
  assign n3415_o = execute_engine[32:28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1097:43  */
  assign n3416_o = execute_engine[39:35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1098:43  */
  assign n3417_o = execute_engine[19:15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1099:31  */
  assign n3418_o = ctrl[22:21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1100:31  */
  assign n3419_o = ctrl[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1103:31  */
  assign n3420_o = ctrl[26:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1104:31  */
  assign n3421_o = ctrl[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1105:31  */
  assign n3422_o = ctrl[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1106:31  */
  assign n3423_o = ctrl[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1107:31  */
  assign n3424_o = ctrl[35:30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1110:31  */
  assign n3425_o = ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1111:31  */
  assign n3426_o = ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1112:51  */
  assign n3428_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1112:57  */
  assign n3430_o = n3428_o == 4'b1011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1112:30  */
  assign n3431_o = n3430_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1113:31  */
  assign n3433_o = ctrl[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1114:30  */
  assign n3434_o = csr[129]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1114:52  */
  assign n3435_o = csr[130]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1114:42  */
  assign n3436_o = n3435_o ? n3434_o : n3437_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1114:81  */
  assign n3437_o = csr[153]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1117:43  */
  assign n3438_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1118:43  */
  assign n3439_o = execute_engine[39:28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1119:43  */
  assign n3440_o = execute_engine[14:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1122:30  */
  assign n3441_o = csr[153]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1124:36  */
  assign n3442_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1125:37  */
  assign n3443_o = debug_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1136:16  */
  assign n3445_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1139:57  */
  assign n3448_o = monitor[19:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1139:66  */
  assign n3450_o = n3448_o + 10'b0000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1144:30  */
  assign n3455_o = monitor[9:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1144:55  */
  assign n3456_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1144:61  */
  assign n3458_o = n3456_o == 4'b0111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1144:34  */
  assign n3459_o = n3458_o ? n3455_o : 10'b0000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1147:29  */
  assign n3461_o = monitor[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1154:14  */
  assign n3463_o = csr[11:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1157:7  */
  assign n3466_o = n3463_o == 12'b100000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1157:26  */
  assign n3468_o = n3463_o == 12'b100000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1157:26  */
  assign n3469_o = n3466_o | n3468_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1157:42  */
  assign n3471_o = n3463_o == 12'b100000000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1157:42  */
  assign n3472_o = n3469_o | n3471_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1157:58  */
  assign n3474_o = n3463_o == 12'b100000000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1157:58  */
  assign n3475_o = n3472_o | n3474_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1161:7  */
  assign n3478_o = n3463_o == 12'b000000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1161:25  */
  assign n3480_o = n3463_o == 12'b000000000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1161:25  */
  assign n3481_o = n3478_o | n3480_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1161:37  */
  assign n3483_o = n3463_o == 12'b000000000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1161:37  */
  assign n3484_o = n3481_o | n3483_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:7  */
  assign n3486_o = n3463_o == 12'b001100000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:27  */
  assign n3488_o = n3463_o == 12'b001100010000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:27  */
  assign n3489_o = n3486_o | n3488_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:49  */
  assign n3491_o = n3463_o == 12'b001100000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:49  */
  assign n3492_o = n3489_o | n3491_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:67  */
  assign n3494_o = n3463_o == 12'b001100000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:67  */
  assign n3495_o = n3492_o | n3494_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:83  */
  assign n3497_o = n3463_o == 12'b001100000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:83  */
  assign n3498_o = n3495_o | n3497_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:98  */
  assign n3500_o = n3463_o == 12'b001101000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1165:98  */
  assign n3501_o = n3498_o | n3500_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:27  */
  assign n3503_o = n3463_o == 12'b001101000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:27  */
  assign n3504_o = n3501_o | n3503_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:49  */
  assign n3506_o = n3463_o == 12'b001101000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:49  */
  assign n3507_o = n3504_o | n3506_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:67  */
  assign n3509_o = n3463_o == 12'b001101000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:67  */
  assign n3510_o = n3507_o | n3509_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:83  */
  assign n3512_o = n3463_o == 12'b001101000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:83  */
  assign n3513_o = n3510_o | n3512_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:98  */
  assign n3515_o = n3463_o == 12'b001101001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1166:98  */
  assign n3516_o = n3513_o | n3515_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:27  */
  assign n3518_o = n3463_o == 12'b001100100000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:27  */
  assign n3519_o = n3516_o | n3518_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:49  */
  assign n3521_o = n3463_o == 12'b111100010001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:49  */
  assign n3522_o = n3519_o | n3521_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:67  */
  assign n3524_o = n3463_o == 12'b111100010010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:67  */
  assign n3525_o = n3522_o | n3524_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:83  */
  assign n3527_o = n3463_o == 12'b111100010011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:83  */
  assign n3528_o = n3525_o | n3527_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:98  */
  assign n3530_o = n3463_o == 12'b111100010100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1167:98  */
  assign n3531_o = n3528_o | n3530_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1168:27  */
  assign n3533_o = n3463_o == 12'b111100010101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1168:27  */
  assign n3534_o = n3531_o | n3533_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1168:49  */
  assign n3536_o = n3463_o == 12'b111111000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1168:49  */
  assign n3537_o = n3534_o | n3536_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1172:7  */
  assign n3540_o = n3463_o == 12'b001100000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1172:29  */
  assign n3542_o = n3463_o == 12'b001100001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1172:29  */
  assign n3543_o = n3540_o | n3542_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1172:45  */
  assign n3545_o = n3463_o == 12'b001100011010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1172:45  */
  assign n3546_o = n3543_o | n3545_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:7  */
  assign n3549_o = n3463_o == 12'b001110100000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:28  */
  assign n3551_o = n3463_o == 12'b001110100001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:28  */
  assign n3552_o = n3549_o | n3551_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:46  */
  assign n3554_o = n3463_o == 12'b001110100010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:46  */
  assign n3555_o = n3552_o | n3554_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:64  */
  assign n3557_o = n3463_o == 12'b001110100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:64  */
  assign n3558_o = n3555_o | n3557_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:82  */
  assign n3560_o = n3463_o == 12'b001110110000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1176:82  */
  assign n3561_o = n3558_o | n3560_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1177:28  */
  assign n3563_o = n3463_o == 12'b001110110001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1177:28  */
  assign n3564_o = n3561_o | n3563_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1177:46  */
  assign n3566_o = n3463_o == 12'b001110110010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1177:46  */
  assign n3567_o = n3564_o | n3566_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1177:64  */
  assign n3569_o = n3463_o == 12'b001110110011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1177:64  */
  assign n3570_o = n3567_o | n3569_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1177:82  */
  assign n3572_o = n3463_o == 12'b001110110100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1177:82  */
  assign n3573_o = n3570_o | n3572_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1178:28  */
  assign n3575_o = n3463_o == 12'b001110110101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1178:28  */
  assign n3576_o = n3573_o | n3575_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1178:46  */
  assign n3578_o = n3463_o == 12'b001110110110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1178:46  */
  assign n3579_o = n3576_o | n3578_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1178:64  */
  assign n3581_o = n3463_o == 12'b001110110111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1178:64  */
  assign n3582_o = n3579_o | n3581_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1178:82  */
  assign n3584_o = n3463_o == 12'b001110111000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1178:82  */
  assign n3585_o = n3582_o | n3584_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1179:28  */
  assign n3587_o = n3463_o == 12'b001110111001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1179:28  */
  assign n3588_o = n3585_o | n3587_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1179:46  */
  assign n3590_o = n3463_o == 12'b001110111010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1179:46  */
  assign n3591_o = n3588_o | n3590_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1179:64  */
  assign n3593_o = n3463_o == 12'b001110111011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1179:64  */
  assign n3594_o = n3591_o | n3593_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1179:82  */
  assign n3596_o = n3463_o == 12'b001110111100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1179:82  */
  assign n3597_o = n3594_o | n3596_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1180:28  */
  assign n3599_o = n3463_o == 12'b001110111101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1180:28  */
  assign n3600_o = n3597_o | n3599_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1180:46  */
  assign n3602_o = n3463_o == 12'b001110111110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1180:46  */
  assign n3603_o = n3600_o | n3602_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1180:64  */
  assign n3605_o = n3463_o == 12'b001110111111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1180:64  */
  assign n3606_o = n3603_o | n3605_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:7  */
  assign n3609_o = n3463_o == 12'b110000000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:33  */
  assign n3611_o = n3463_o == 12'b110000000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:33  */
  assign n3612_o = n3609_o | n3611_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:56  */
  assign n3614_o = n3463_o == 12'b110000000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:56  */
  assign n3615_o = n3612_o | n3614_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:79  */
  assign n3617_o = n3463_o == 12'b110000000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:79  */
  assign n3618_o = n3615_o | n3617_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:102  */
  assign n3620_o = n3463_o == 12'b110000000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:102  */
  assign n3621_o = n3618_o | n3620_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:125  */
  assign n3623_o = n3463_o == 12'b110000001000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1184:125  */
  assign n3624_o = n3621_o | n3623_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:33  */
  assign n3626_o = n3463_o == 12'b110000001001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:33  */
  assign n3627_o = n3624_o | n3626_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:56  */
  assign n3629_o = n3463_o == 12'b110000001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:56  */
  assign n3630_o = n3627_o | n3629_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:79  */
  assign n3632_o = n3463_o == 12'b110000001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:79  */
  assign n3633_o = n3630_o | n3632_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:102  */
  assign n3635_o = n3463_o == 12'b110000001100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:102  */
  assign n3636_o = n3633_o | n3635_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:125  */
  assign n3638_o = n3463_o == 12'b110000001101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1185:125  */
  assign n3639_o = n3636_o | n3638_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1186:33  */
  assign n3641_o = n3463_o == 12'b110000001110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1186:33  */
  assign n3642_o = n3639_o | n3641_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1186:56  */
  assign n3644_o = n3463_o == 12'b110000001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1186:56  */
  assign n3645_o = n3642_o | n3644_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1186:79  */
  assign n3647_o = n3463_o == 12'b110010000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1186:79  */
  assign n3648_o = n3645_o | n3647_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:33  */
  assign n3650_o = n3463_o == 12'b110010000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:33  */
  assign n3651_o = n3648_o | n3650_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:56  */
  assign n3653_o = n3463_o == 12'b110010000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:56  */
  assign n3654_o = n3651_o | n3653_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:79  */
  assign n3656_o = n3463_o == 12'b110010000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:79  */
  assign n3657_o = n3654_o | n3656_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:102  */
  assign n3659_o = n3463_o == 12'b110010000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:102  */
  assign n3660_o = n3657_o | n3659_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:125  */
  assign n3662_o = n3463_o == 12'b110010001000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1187:125  */
  assign n3663_o = n3660_o | n3662_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:33  */
  assign n3665_o = n3463_o == 12'b110010001001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:33  */
  assign n3666_o = n3663_o | n3665_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:56  */
  assign n3668_o = n3463_o == 12'b110010001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:56  */
  assign n3669_o = n3666_o | n3668_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:79  */
  assign n3671_o = n3463_o == 12'b110010001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:79  */
  assign n3672_o = n3669_o | n3671_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:102  */
  assign n3674_o = n3463_o == 12'b110010001100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:102  */
  assign n3675_o = n3672_o | n3674_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:125  */
  assign n3677_o = n3463_o == 12'b110010001101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1188:125  */
  assign n3678_o = n3675_o | n3677_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1189:33  */
  assign n3680_o = n3463_o == 12'b110010001110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1189:33  */
  assign n3681_o = n3678_o | n3680_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1189:56  */
  assign n3683_o = n3463_o == 12'b110010001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1189:56  */
  assign n3684_o = n3681_o | n3683_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1189:79  */
  assign n3686_o = n3463_o == 12'b101100000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1189:79  */
  assign n3687_o = n3684_o | n3686_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:33  */
  assign n3689_o = n3463_o == 12'b101100000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:33  */
  assign n3690_o = n3687_o | n3689_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:56  */
  assign n3692_o = n3463_o == 12'b101100000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:56  */
  assign n3693_o = n3690_o | n3692_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:79  */
  assign n3695_o = n3463_o == 12'b101100000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:79  */
  assign n3696_o = n3693_o | n3695_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:102  */
  assign n3698_o = n3463_o == 12'b101100000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:102  */
  assign n3699_o = n3696_o | n3698_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:125  */
  assign n3701_o = n3463_o == 12'b101100001000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1190:125  */
  assign n3702_o = n3699_o | n3701_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:33  */
  assign n3704_o = n3463_o == 12'b101100001001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:33  */
  assign n3705_o = n3702_o | n3704_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:56  */
  assign n3707_o = n3463_o == 12'b101100001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:56  */
  assign n3708_o = n3705_o | n3707_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:79  */
  assign n3710_o = n3463_o == 12'b101100001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:79  */
  assign n3711_o = n3708_o | n3710_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:102  */
  assign n3713_o = n3463_o == 12'b101100001100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:102  */
  assign n3714_o = n3711_o | n3713_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:125  */
  assign n3716_o = n3463_o == 12'b101100001101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1191:125  */
  assign n3717_o = n3714_o | n3716_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1192:33  */
  assign n3719_o = n3463_o == 12'b101100001110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1192:33  */
  assign n3720_o = n3717_o | n3719_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1192:56  */
  assign n3722_o = n3463_o == 12'b101100001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1192:56  */
  assign n3723_o = n3720_o | n3722_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1192:79  */
  assign n3725_o = n3463_o == 12'b101110000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1192:79  */
  assign n3726_o = n3723_o | n3725_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:33  */
  assign n3728_o = n3463_o == 12'b101110000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:33  */
  assign n3729_o = n3726_o | n3728_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:56  */
  assign n3731_o = n3463_o == 12'b101110000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:56  */
  assign n3732_o = n3729_o | n3731_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:79  */
  assign n3734_o = n3463_o == 12'b101110000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:79  */
  assign n3735_o = n3732_o | n3734_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:102  */
  assign n3737_o = n3463_o == 12'b101110000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:102  */
  assign n3738_o = n3735_o | n3737_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:125  */
  assign n3740_o = n3463_o == 12'b101110001000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1193:125  */
  assign n3741_o = n3738_o | n3740_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:33  */
  assign n3743_o = n3463_o == 12'b101110001001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:33  */
  assign n3744_o = n3741_o | n3743_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:56  */
  assign n3746_o = n3463_o == 12'b101110001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:56  */
  assign n3747_o = n3744_o | n3746_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:79  */
  assign n3749_o = n3463_o == 12'b101110001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:79  */
  assign n3750_o = n3747_o | n3749_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:102  */
  assign n3752_o = n3463_o == 12'b101110001100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:102  */
  assign n3753_o = n3750_o | n3752_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:125  */
  assign n3755_o = n3463_o == 12'b101110001101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1194:125  */
  assign n3756_o = n3753_o | n3755_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1195:33  */
  assign n3758_o = n3463_o == 12'b101110001110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1195:33  */
  assign n3759_o = n3756_o | n3758_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1195:56  */
  assign n3761_o = n3463_o == 12'b101110001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1195:56  */
  assign n3762_o = n3759_o | n3761_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1195:79  */
  assign n3764_o = n3463_o == 12'b001100100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1195:79  */
  assign n3765_o = n3762_o | n3764_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:33  */
  assign n3767_o = n3463_o == 12'b001100100100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:33  */
  assign n3768_o = n3765_o | n3767_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:56  */
  assign n3770_o = n3463_o == 12'b001100100101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:56  */
  assign n3771_o = n3768_o | n3770_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:79  */
  assign n3773_o = n3463_o == 12'b001100100110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:79  */
  assign n3774_o = n3771_o | n3773_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:102  */
  assign n3776_o = n3463_o == 12'b001100100111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:102  */
  assign n3777_o = n3774_o | n3776_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:125  */
  assign n3779_o = n3463_o == 12'b001100101000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1196:125  */
  assign n3780_o = n3777_o | n3779_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:33  */
  assign n3782_o = n3463_o == 12'b001100101001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:33  */
  assign n3783_o = n3780_o | n3782_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:56  */
  assign n3785_o = n3463_o == 12'b001100101010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:56  */
  assign n3786_o = n3783_o | n3785_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:79  */
  assign n3788_o = n3463_o == 12'b001100101011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:79  */
  assign n3789_o = n3786_o | n3788_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:102  */
  assign n3791_o = n3463_o == 12'b001100101100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:102  */
  assign n3792_o = n3789_o | n3791_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:125  */
  assign n3794_o = n3463_o == 12'b001100101101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1197:125  */
  assign n3795_o = n3792_o | n3794_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1198:33  */
  assign n3797_o = n3463_o == 12'b001100101110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1198:33  */
  assign n3798_o = n3795_o | n3797_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1198:56  */
  assign n3800_o = n3463_o == 12'b001100101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1198:56  */
  assign n3801_o = n3798_o | n3800_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:7  */
  assign n3804_o = n3463_o == 12'b110000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:25  */
  assign n3806_o = n3463_o == 12'b101100000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:25  */
  assign n3807_o = n3804_o | n3806_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:41  */
  assign n3809_o = n3463_o == 12'b110000000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:41  */
  assign n3810_o = n3807_o | n3809_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:58  */
  assign n3812_o = n3463_o == 12'b101100000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:58  */
  assign n3813_o = n3810_o | n3812_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:75  */
  assign n3815_o = n3463_o == 12'b110010000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1202:75  */
  assign n3816_o = n3813_o | n3815_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1203:25  */
  assign n3818_o = n3463_o == 12'b101110000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1203:25  */
  assign n3819_o = n3816_o | n3818_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1203:41  */
  assign n3821_o = n3463_o == 12'b110010000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1203:41  */
  assign n3822_o = n3819_o | n3821_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1203:58  */
  assign n3824_o = n3463_o == 12'b101110000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1203:58  */
  assign n3825_o = n3822_o | n3824_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1207:7  */
  assign n3828_o = n3463_o == 12'b011110110000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1207:23  */
  assign n3830_o = n3463_o == 12'b011110110001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1207:23  */
  assign n3831_o = n3828_o | n3830_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1207:35  */
  assign n3833_o = n3463_o == 12'b011110110010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1207:35  */
  assign n3834_o = n3831_o | n3833_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1211:7  */
  assign n3837_o = n3463_o == 12'b011110100000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1211:26  */
  assign n3839_o = n3463_o == 12'b011110100001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1211:26  */
  assign n3840_o = n3837_o | n3839_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1211:41  */
  assign n3842_o = n3463_o == 12'b011110100010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1211:41  */
  assign n3843_o = n3840_o | n3842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1211:56  */
  assign n3845_o = n3463_o == 12'b011110100100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1211:56  */
  assign n3846_o = n3843_o | n3845_o;
  assign n3847_o = {n3846_o, n3834_o, n3825_o, n3801_o, n3606_o, n3546_o, n3537_o, n3484_o, n3475_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1154:5  */
  always @*
    case (n3847_o)
      9'b100000000: n3858_o = 1'b0;
      9'b010000000: n3858_o = 1'b0;
      9'b001000000: n3858_o = 1'b1;
      9'b000100000: n3858_o = 1'b0;
      9'b000010000: n3858_o = 1'b0;
      9'b000001000: n3858_o = 1'b1;
      9'b000000100: n3858_o = 1'b1;
      9'b000000010: n3858_o = 1'b0;
      9'b000000001: n3858_o = 1'b0;
      default: n3858_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1226:17  */
  assign n3861_o = csr[11:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1226:32  */
  assign n3863_o = n3861_o == 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1227:27  */
  assign n3864_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1227:74  */
  assign n3866_o = n3864_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1228:27  */
  assign n3867_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1228:74  */
  assign n3869_o = n3867_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1227:93  */
  assign n3870_o = n3866_o | n3869_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1229:21  */
  assign n3871_o = decode_aux[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1229:30  */
  assign n3872_o = ~n3871_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1228:93  */
  assign n3873_o = n3870_o | n3872_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1226:40  */
  assign n3874_o = n3873_o & n3863_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1226:5  */
  assign n3877_o = n3874_o ? 1'b0 : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1244:20  */
  assign n3891_o = csr[11:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1244:34  */
  assign n3893_o = n3891_o == 4'b1100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1244:62  */
  assign n3895_o = 1'b1 & n3893_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1245:87  */
  assign n3897_o = 1'b1 & n3895_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1246:51  */
  assign n3898_o = csr[153]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1246:65  */
  assign n3899_o = ~n3898_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1246:42  */
  assign n3900_o = n3899_o & n3897_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1246:81  */
  assign n3901_o = csr[320]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1246:92  */
  assign n3902_o = ~n3901_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1246:72  */
  assign n3903_o = n3902_o & n3900_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1248:20  */
  assign n3904_o = csr[9:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1248:33  */
  assign n3906_o = n3904_o != 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1248:51  */
  assign n3907_o = csr[153]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1248:65  */
  assign n3908_o = ~n3907_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1248:42  */
  assign n3909_o = n3908_o & n3906_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1248:5  */
  assign n3912_o = n3909_o ? 1'b0 : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1244:5  */
  assign n3914_o = n3903_o ? 1'b0 : n3912_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1261:21  */
  assign n3917_o = decode_aux[6:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1263:7  */
  assign n3919_o = n3917_o == 7'b0110111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1263:25  */
  assign n3921_o = n3917_o == 7'b0010111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1263:25  */
  assign n3922_o = n3919_o | n3921_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1263:42  */
  assign n3924_o = n3917_o == 7'b1101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1263:42  */
  assign n3925_o = n3922_o | n3924_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1267:31  */
  assign n3926_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1268:11  */
  assign n3928_o = n3926_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1267:9  */
  always @*
    case (n3928_o)
      1'b1: n3931_o = 1'b0;
      default: n3931_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1266:7  */
  assign n3933_o = n3917_o == 7'b1100111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1273:31  */
  assign n3934_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:11  */
  assign n3936_o = n3934_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:29  */
  assign n3938_o = n3934_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:29  */
  assign n3939_o = n3936_o | n3938_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:44  */
  assign n3941_o = n3934_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:44  */
  assign n3942_o = n3939_o | n3941_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:59  */
  assign n3944_o = n3934_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:59  */
  assign n3945_o = n3942_o | n3944_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:74  */
  assign n3947_o = n3934_o == 3'b110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:74  */
  assign n3948_o = n3945_o | n3947_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:90  */
  assign n3950_o = n3934_o == 3'b111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1274:90  */
  assign n3951_o = n3948_o | n3950_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1273:9  */
  always @*
    case (n3951_o)
      1'b1: n3954_o = 1'b0;
      default: n3954_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1272:7  */
  assign n3956_o = n3917_o == 7'b1100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1279:31  */
  assign n3957_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:11  */
  assign n3959_o = n3957_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:28  */
  assign n3961_o = n3957_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:28  */
  assign n3962_o = n3959_o | n3961_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:42  */
  assign n3964_o = n3957_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:42  */
  assign n3965_o = n3962_o | n3964_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:56  */
  assign n3967_o = n3957_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:56  */
  assign n3968_o = n3965_o | n3967_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:71  */
  assign n3970_o = n3957_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1280:71  */
  assign n3971_o = n3968_o | n3970_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1279:9  */
  always @*
    case (n3971_o)
      1'b1: n3974_o = 1'b0;
      default: n3974_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1278:7  */
  assign n3976_o = n3917_o == 7'b0000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1285:31  */
  assign n3977_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1286:11  */
  assign n3979_o = n3977_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1286:28  */
  assign n3981_o = n3977_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1286:28  */
  assign n3982_o = n3979_o | n3981_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1286:42  */
  assign n3984_o = n3977_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1286:42  */
  assign n3985_o = n3982_o | n3984_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1285:9  */
  always @*
    case (n3985_o)
      1'b1: n3988_o = 1'b0;
      default: n3988_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1284:7  */
  assign n3990_o = n3917_o == 7'b0100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1290:7  */
  assign n3992_o = n3917_o == 7'b0101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1298:33  */
  assign n3993_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1298:80  */
  assign n3995_o = n3993_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1298:120  */
  assign n3996_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1298:167  */
  assign n3998_o = n3996_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1298:99  */
  assign n3999_o = n3995_o | n3998_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1299:32  */
  assign n4000_o = execute_engine[37:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1299:81  */
  assign n4002_o = n4000_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1298:183  */
  assign n4003_o = n4002_o & n3999_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1299:114  */
  assign n4004_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1299:135  */
  assign n4005_o = ~n4004_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1299:92  */
  assign n4006_o = n4005_o & n4003_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1300:33  */
  assign n4007_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1300:80  */
  assign n4009_o = n4007_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1301:33  */
  assign n4010_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1301:80  */
  assign n4012_o = n4010_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1300:96  */
  assign n4013_o = n4009_o | n4012_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1302:33  */
  assign n4014_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1302:80  */
  assign n4016_o = n4014_o == 3'b011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1301:96  */
  assign n4017_o = n4013_o | n4016_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1303:33  */
  assign n4018_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1303:80  */
  assign n4020_o = n4018_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1302:97  */
  assign n4021_o = n4017_o | n4020_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1304:33  */
  assign n4022_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1304:80  */
  assign n4024_o = n4022_o == 3'b110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1303:96  */
  assign n4025_o = n4021_o | n4024_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1305:33  */
  assign n4026_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1305:80  */
  assign n4028_o = n4026_o == 3'b111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1304:95  */
  assign n4029_o = n4025_o | n4028_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1306:33  */
  assign n4030_o = execute_engine[39:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1306:80  */
  assign n4032_o = n4030_o == 7'b0000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1305:97  */
  assign n4033_o = n4032_o & n4029_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1299:143  */
  assign n4034_o = n4006_o | n4033_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1307:100  */
  assign n4035_o = decode_aux[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1307:84  */
  assign n4037_o = n4035_o & 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1306:95  */
  assign n4038_o = n4034_o | n4037_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1308:60  */
  assign n4039_o = decode_aux[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1308:44  */
  assign n4041_o = n4039_o & 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1307:117  */
  assign n4042_o = n4038_o | n4041_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1308:77  */
  assign n4044_o = n4042_o | 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1309:77  */
  assign n4046_o = n4044_o | 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1298:9  */
  assign n4049_o = n4046_o ? 1'b0 : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1297:7  */
  assign n4051_o = n3917_o == 7'b0110011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1317:31  */
  assign n4052_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1317:78  */
  assign n4054_o = n4052_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1318:31  */
  assign n4055_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1318:78  */
  assign n4057_o = n4055_o == 3'b010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1317:97  */
  assign n4058_o = n4054_o | n4057_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1319:31  */
  assign n4059_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1319:78  */
  assign n4061_o = n4059_o == 3'b011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1318:94  */
  assign n4062_o = n4058_o | n4061_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1320:31  */
  assign n4063_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1320:78  */
  assign n4065_o = n4063_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1319:95  */
  assign n4066_o = n4062_o | n4065_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1321:31  */
  assign n4067_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1321:78  */
  assign n4069_o = n4067_o == 3'b110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1320:94  */
  assign n4070_o = n4066_o | n4069_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1322:31  */
  assign n4071_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1322:78  */
  assign n4073_o = n4071_o == 3'b111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1321:93  */
  assign n4074_o = n4070_o | n4073_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1323:32  */
  assign n4075_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1323:79  */
  assign n4077_o = n4075_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1324:32  */
  assign n4078_o = execute_engine[39:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1324:79  */
  assign n4080_o = n4078_o == 7'b0000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1323:95  */
  assign n4081_o = n4080_o & n4077_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1322:94  */
  assign n4082_o = n4074_o | n4081_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1325:32  */
  assign n4083_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1325:79  */
  assign n4085_o = n4083_o == 3'b101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1326:33  */
  assign n4086_o = execute_engine[37:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1326:82  */
  assign n4088_o = n4086_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1326:115  */
  assign n4089_o = execute_engine[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1326:136  */
  assign n4090_o = ~n4089_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1326:93  */
  assign n4091_o = n4090_o & n4088_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1325:94  */
  assign n4092_o = n4091_o & n4085_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1324:93  */
  assign n4093_o = n4082_o | n4092_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1326:146  */
  assign n4095_o = n4093_o | 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1317:9  */
  assign n4098_o = n4095_o ? 1'b0 : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1316:7  */
  assign n4100_o = n3917_o == 7'b0010011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1334:31  */
  assign n4101_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1335:11  */
  assign n4103_o = n4101_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1335:31  */
  assign n4105_o = n4101_o == 3'b001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1335:31  */
  assign n4106_o = n4103_o | n4105_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1334:9  */
  always @*
    case (n4106_o)
      1'b1: n4109_o = 1'b0;
      default: n4109_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1333:7  */
  assign n4111_o = n3917_o == 7'b0001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1340:30  */
  assign n4112_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1340:77  */
  assign n4114_o = n4112_o == 3'b000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1341:26  */
  assign n4115_o = decode_aux[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1341:58  */
  assign n4116_o = decode_aux[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1341:42  */
  assign n4117_o = n4116_o & n4115_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1342:35  */
  assign n4118_o = execute_engine[39:28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1343:15  */
  assign n4120_o = n4118_o == 12'b000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1343:36  */
  assign n4122_o = n4118_o == 12'b000000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1343:36  */
  assign n4123_o = n4120_o | n4122_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1344:82  */
  assign n4124_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1344:74  */
  assign n4125_o = ~n4124_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1344:107  */
  assign n4126_o = debug_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1344:93  */
  assign n4127_o = n4125_o | n4126_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1344:15  */
  assign n4129_o = n4118_o == 12'b001100000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1345:88  */
  assign n4130_o = debug_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1345:73  */
  assign n4131_o = ~n4130_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1345:15  */
  assign n4133_o = n4118_o == 12'b011110110010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1346:82  */
  assign n4134_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1346:74  */
  assign n4135_o = ~n4134_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1346:101  */
  assign n4136_o = csr[131]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1346:93  */
  assign n4137_o = n4135_o & n4136_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1346:15  */
  assign n4139_o = n4118_o == 12'b000100000101;
  assign n4140_o = {n4139_o, n4133_o, n4129_o, n4123_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1342:13  */
  always @*
    case (n4140_o)
      4'b1000: n4143_o = n4137_o;
      4'b0100: n4143_o = n4131_o;
      4'b0010: n4143_o = n4127_o;
      4'b0001: n4143_o = 1'b0;
      default: n4143_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1341:11  */
  assign n4145_o = n4117_o ? n4143_o : 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1352:30  */
  assign n4146_o = ~csr_reg_valid;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1352:54  */
  assign n4147_o = ~csr_rw_valid;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1352:37  */
  assign n4148_o = n4146_o | n4147_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1352:80  */
  assign n4149_o = ~csr_priv_valid;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1352:61  */
  assign n4150_o = n4148_o | n4149_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1353:33  */
  assign n4151_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1353:80  */
  assign n4153_o = n4151_o == 3'b100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1352:87  */
  assign n4154_o = n4150_o | n4153_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1352:9  */
  assign n4157_o = n4154_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1340:9  */
  assign n4158_o = n4114_o ? n4145_o : n4157_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1339:7  */
  assign n4160_o = n3917_o == 7'b1110011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1360:93  */
  assign n4162_o = decode_aux[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1360:78  */
  assign n4163_o = ~n4162_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1360:74  */
  assign n4165_o = 1'b1 | n4163_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1359:7  */
  assign n4167_o = n3917_o == 7'b1010011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1362:7  */
  assign n4170_o = n3917_o == 7'b0001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1362:27  */
  assign n4172_o = n3917_o == 7'b0101011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1362:27  */
  assign n4173_o = n4170_o | n4172_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1362:44  */
  assign n4175_o = n3917_o == 7'b1011011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1362:44  */
  assign n4176_o = n4173_o | n4175_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1362:61  */
  assign n4178_o = n3917_o == 7'b1111011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1362:61  */
  assign n4179_o = n4176_o | n4178_o;
  assign n4180_o = {n4179_o, n4167_o, n4160_o, n4111_o, n4100_o, n4051_o, n3992_o, n3990_o, n3976_o, n3956_o, n3933_o, n3925_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1261:5  */
  always @*
    case (n4180_o)
      12'b100000000000: n4185_o = 1'b1;
      12'b010000000000: n4185_o = n4165_o;
      12'b001000000000: n4185_o = n4158_o;
      12'b000100000000: n4185_o = n4109_o;
      12'b000010000000: n4185_o = n4098_o;
      12'b000001000000: n4185_o = n4049_o;
      12'b000000100000: n4185_o = 1'b1;
      12'b000000010000: n4185_o = n3988_o;
      12'b000000001000: n4185_o = n3974_o;
      12'b000000000100: n4185_o = n3954_o;
      12'b000000000010: n4185_o = n3931_o;
      12'b000000000001: n4185_o = 1'b0;
      default: n4185_o = 1'b1;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1374:51  */
  assign n4189_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1374:57  */
  assign n4191_o = n4189_o == 4'b0110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1374:87  */
  assign n4192_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1374:93  */
  assign n4194_o = n4192_o == 4'b0111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1374:68  */
  assign n4195_o = n4191_o | n4194_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1375:44  */
  assign n4196_o = monitor[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1375:55  */
  assign n4197_o = n4196_o | illegal_cmd;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1377:53  */
  assign n4198_o = execute_engine[9:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1377:102  */
  assign n4200_o = n4198_o != 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1376:55  */
  assign n4201_o = n4197_o | n4200_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1374:106  */
  assign n4202_o = n4201_o & n4195_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1374:29  */
  assign n4203_o = n4202_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1388:16  */
  assign n4206_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1400:60  */
  assign n4209_o = trap_ctrl[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1400:75  */
  assign n4210_o = n4209_o | ma_load_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1400:117  */
  assign n4211_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1400:103  */
  assign n4212_o = ~n4211_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1400:98  */
  assign n4213_o = n4210_o & n4212_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1401:60  */
  assign n4214_o = trap_ctrl[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1401:75  */
  assign n4215_o = n4214_o | ma_store_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1401:117  */
  assign n4216_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1401:103  */
  assign n4217_o = ~n4216_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1401:98  */
  assign n4218_o = n4215_o & n4217_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1402:60  */
  assign n4219_o = trap_ctrl[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1402:88  */
  assign n4220_o = trap_ctrl[99]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1402:75  */
  assign n4221_o = n4219_o | n4220_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1402:117  */
  assign n4222_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1402:103  */
  assign n4223_o = ~n4222_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1402:98  */
  assign n4224_o = n4221_o & n4223_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1405:61  */
  assign n4225_o = trap_ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1405:77  */
  assign n4226_o = n4225_o | be_load_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1405:119  */
  assign n4227_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1405:105  */
  assign n4228_o = ~n4227_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1405:100  */
  assign n4229_o = n4226_o & n4228_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1406:61  */
  assign n4230_o = trap_ctrl[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1406:77  */
  assign n4231_o = n4230_o | be_store_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1406:119  */
  assign n4232_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1406:105  */
  assign n4233_o = ~n4232_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1406:100  */
  assign n4234_o = n4231_o & n4233_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1407:61  */
  assign n4235_o = trap_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1407:90  */
  assign n4236_o = trap_ctrl[98]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1407:77  */
  assign n4237_o = n4235_o | n4236_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1407:119  */
  assign n4238_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1407:105  */
  assign n4239_o = ~n4238_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1407:100  */
  assign n4240_o = n4237_o & n4239_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1410:61  */
  assign n4241_o = trap_ctrl[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1410:90  */
  assign n4242_o = trap_ctrl[101]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1410:77  */
  assign n4243_o = n4241_o | n4242_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1410:119  */
  assign n4244_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1410:105  */
  assign n4245_o = ~n4244_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1410:100  */
  assign n4246_o = n4243_o & n4245_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1411:61  */
  assign n4247_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1411:90  */
  assign n4248_o = trap_ctrl[100]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1411:77  */
  assign n4249_o = n4247_o | n4248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1411:119  */
  assign n4250_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1411:105  */
  assign n4251_o = ~n4250_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1411:100  */
  assign n4252_o = n4249_o & n4251_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:62  */
  assign n4253_o = trap_ctrl[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:90  */
  assign n4254_o = trap_ctrl[102]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:77  */
  assign n4255_o = n4253_o | n4254_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:111  */
  assign n4256_o = trap_ctrl[103]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:131  */
  assign n4257_o = csr[442]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:123  */
  assign n4258_o = ~n4257_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:118  */
  assign n4259_o = n4256_o & n4258_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:97  */
  assign n4260_o = n4255_o | n4259_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:167  */
  assign n4261_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:153  */
  assign n4262_o = ~n4261_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1420:148  */
  assign n4263_o = n4260_o & n4262_o;
  assign n4266_o = {1'b0, 1'b0, n4229_o, n4234_o, n4213_o, n4218_o, n4263_o, n4246_o, n4224_o, n4252_o, n4240_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1439:16  */
  assign n4272_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4276_o = firq_i[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4278_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4279_o = csr[111]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4280_o = ~n4279_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4281_o = n4280_o & n4278_o;
  assign n4283_o = trap_ctrl[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4284_o = n4281_o ? 1'b0 : n4283_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4285_o = n4276_o ? 1'b1 : n4284_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4286_o = firq_i[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4288_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4289_o = csr[112]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4290_o = ~n4289_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4291_o = n4290_o & n4288_o;
  assign n4293_o = trap_ctrl[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4294_o = n4291_o ? 1'b0 : n4293_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4295_o = n4286_o ? 1'b1 : n4294_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4296_o = firq_i[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4298_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4299_o = csr[113]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4300_o = ~n4299_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4301_o = n4300_o & n4298_o;
  assign n4303_o = trap_ctrl[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4304_o = n4301_o ? 1'b0 : n4303_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4305_o = n4296_o ? 1'b1 : n4304_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4306_o = firq_i[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4308_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4309_o = csr[114]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4310_o = ~n4309_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4311_o = n4310_o & n4308_o;
  assign n4313_o = trap_ctrl[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4314_o = n4311_o ? 1'b0 : n4313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4315_o = n4306_o ? 1'b1 : n4314_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4316_o = firq_i[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4318_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4319_o = csr[115]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4320_o = ~n4319_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4321_o = n4320_o & n4318_o;
  assign n4323_o = trap_ctrl[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4324_o = n4321_o ? 1'b0 : n4323_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4325_o = n4316_o ? 1'b1 : n4324_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4326_o = firq_i[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4328_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4329_o = csr[116]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4330_o = ~n4329_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4331_o = n4330_o & n4328_o;
  assign n4333_o = trap_ctrl[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4334_o = n4331_o ? 1'b0 : n4333_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4335_o = n4326_o ? 1'b1 : n4334_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4336_o = firq_i[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4338_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4339_o = csr[117]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4340_o = ~n4339_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4341_o = n4340_o & n4338_o;
  assign n4343_o = trap_ctrl[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4344_o = n4341_o ? 1'b0 : n4343_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4345_o = n4336_o ? 1'b1 : n4344_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4346_o = firq_i[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4348_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4349_o = csr[118]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4350_o = ~n4349_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4351_o = n4350_o & n4348_o;
  assign n4353_o = trap_ctrl[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4354_o = n4351_o ? 1'b0 : n4353_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4355_o = n4346_o ? 1'b1 : n4354_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4356_o = firq_i[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4358_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4359_o = csr[119]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4360_o = ~n4359_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4361_o = n4360_o & n4358_o;
  assign n4363_o = trap_ctrl[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4364_o = n4361_o ? 1'b0 : n4363_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4365_o = n4356_o ? 1'b1 : n4364_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4366_o = firq_i[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4368_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4369_o = csr[120]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4370_o = ~n4369_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4371_o = n4370_o & n4368_o;
  assign n4373_o = trap_ctrl[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4374_o = n4371_o ? 1'b0 : n4373_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4375_o = n4366_o ? 1'b1 : n4374_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4376_o = firq_i[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4378_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4379_o = csr[121]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4380_o = ~n4379_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4381_o = n4380_o & n4378_o;
  assign n4383_o = trap_ctrl[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4384_o = n4381_o ? 1'b0 : n4383_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4385_o = n4376_o ? 1'b1 : n4384_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4386_o = firq_i[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4388_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4389_o = csr[122]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4390_o = ~n4389_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4391_o = n4390_o & n4388_o;
  assign n4393_o = trap_ctrl[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4394_o = n4391_o ? 1'b0 : n4393_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4395_o = n4386_o ? 1'b1 : n4394_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4396_o = firq_i[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4398_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4399_o = csr[123]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4400_o = ~n4399_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4401_o = n4400_o & n4398_o;
  assign n4403_o = trap_ctrl[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4404_o = n4401_o ? 1'b0 : n4403_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4405_o = n4396_o ? 1'b1 : n4404_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4406_o = firq_i[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4408_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4409_o = csr[124]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4410_o = ~n4409_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4411_o = n4410_o & n4408_o;
  assign n4413_o = trap_ctrl[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4414_o = n4411_o ? 1'b0 : n4413_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4415_o = n4406_o ? 1'b1 : n4414_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4416_o = firq_i[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4418_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4419_o = csr[125]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4420_o = ~n4419_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4421_o = n4420_o & n4418_o;
  assign n4423_o = trap_ctrl[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4424_o = n4421_o ? 1'b0 : n4423_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4425_o = n4416_o ? 1'b1 : n4424_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:19  */
  assign n4426_o = firq_i[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:20  */
  assign n4428_o = csr[151]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:53  */
  assign n4429_o = csr[126]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:60  */
  assign n4430_o = ~n4429_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:39  */
  assign n4431_o = n4430_o & n4428_o;
  assign n4433_o = trap_ctrl[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1459:9  */
  assign n4434_o = n4431_o ? 1'b0 : n4433_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1457:9  */
  assign n4435_o = n4426_o ? 1'b1 : n4434_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1475:61  */
  assign n4438_o = trap_ctrl[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1475:85  */
  assign n4439_o = csr[132]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1475:77  */
  assign n4440_o = n4438_o & n4439_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1475:108  */
  assign n4441_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1475:141  */
  assign n4442_o = trap_ctrl[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1475:120  */
  assign n4443_o = n4441_o & n4442_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1475:94  */
  assign n4444_o = n4440_o | n4443_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1476:61  */
  assign n4445_o = trap_ctrl[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1476:85  */
  assign n4446_o = csr[133]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1476:77  */
  assign n4447_o = n4445_o & n4446_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1476:108  */
  assign n4448_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1476:141  */
  assign n4449_o = trap_ctrl[35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1476:120  */
  assign n4450_o = n4448_o & n4449_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1476:94  */
  assign n4451_o = n4447_o | n4450_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1477:61  */
  assign n4452_o = trap_ctrl[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1477:85  */
  assign n4453_o = csr[134]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1477:77  */
  assign n4454_o = n4452_o & n4453_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1477:108  */
  assign n4455_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1477:141  */
  assign n4456_o = trap_ctrl[34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1477:120  */
  assign n4457_o = n4455_o & n4456_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1477:94  */
  assign n4458_o = n4454_o | n4457_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4459_o = trap_ctrl[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4460_o = csr[135]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4461_o = n4459_o & n4460_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4462_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4463_o = trap_ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4464_o = n4462_o & n4463_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4465_o = n4461_o | n4464_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4466_o = trap_ctrl[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4467_o = csr[136]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4468_o = n4466_o & n4467_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4469_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4470_o = trap_ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4471_o = n4469_o & n4470_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4472_o = n4468_o | n4471_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4473_o = trap_ctrl[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4474_o = csr[137]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4475_o = n4473_o & n4474_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4476_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4477_o = trap_ctrl[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4478_o = n4476_o & n4477_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4479_o = n4475_o | n4478_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4480_o = trap_ctrl[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4481_o = csr[138]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4482_o = n4480_o & n4481_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4483_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4484_o = trap_ctrl[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4485_o = n4483_o & n4484_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4486_o = n4482_o | n4485_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4487_o = trap_ctrl[19]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4488_o = csr[139]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4489_o = n4487_o & n4488_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4490_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4491_o = trap_ctrl[40]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4492_o = n4490_o & n4491_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4493_o = n4489_o | n4492_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4494_o = trap_ctrl[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4495_o = csr[140]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4496_o = n4494_o & n4495_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4497_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4498_o = trap_ctrl[41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4499_o = n4497_o & n4498_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4500_o = n4496_o | n4499_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4501_o = trap_ctrl[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4502_o = csr[141]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4503_o = n4501_o & n4502_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4504_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4505_o = trap_ctrl[42]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4506_o = n4504_o & n4505_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4507_o = n4503_o | n4506_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4508_o = trap_ctrl[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4509_o = csr[142]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4510_o = n4508_o & n4509_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4511_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4512_o = trap_ctrl[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4513_o = n4511_o & n4512_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4514_o = n4510_o | n4513_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4515_o = trap_ctrl[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4516_o = csr[143]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4517_o = n4515_o & n4516_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4518_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4519_o = trap_ctrl[44]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4520_o = n4518_o & n4519_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4521_o = n4517_o | n4520_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4522_o = trap_ctrl[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4523_o = csr[144]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4524_o = n4522_o & n4523_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4525_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4526_o = trap_ctrl[45]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4527_o = n4525_o & n4526_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4528_o = n4524_o | n4527_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4529_o = trap_ctrl[25]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4530_o = csr[145]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4531_o = n4529_o & n4530_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4532_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4533_o = trap_ctrl[46]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4534_o = n4532_o & n4533_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4535_o = n4531_o | n4534_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4536_o = trap_ctrl[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4537_o = csr[146]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4538_o = n4536_o & n4537_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4539_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4540_o = trap_ctrl[47]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4541_o = n4539_o & n4540_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4542_o = n4538_o | n4541_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4543_o = trap_ctrl[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4544_o = csr[147]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4545_o = n4543_o & n4544_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4546_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4547_o = trap_ctrl[48]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4548_o = n4546_o & n4547_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4549_o = n4545_o | n4548_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4550_o = trap_ctrl[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4551_o = csr[148]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4552_o = n4550_o & n4551_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4553_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4554_o = trap_ctrl[49]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4555_o = n4553_o & n4554_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4556_o = n4552_o | n4555_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4557_o = trap_ctrl[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4558_o = csr[149]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4559_o = n4557_o & n4558_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4560_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4561_o = trap_ctrl[50]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4562_o = n4560_o & n4561_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4563_o = n4559_o | n4562_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:64  */
  assign n4564_o = trap_ctrl[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:97  */
  assign n4565_o = csr[150]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:81  */
  assign n4566_o = n4564_o & n4565_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:116  */
  assign n4567_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:149  */
  assign n4568_o = trap_ctrl[51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:128  */
  assign n4569_o = n4567_o & n4568_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1481:102  */
  assign n4570_o = n4566_o | n4569_o;
  assign n4573_o = {1'b0, 1'b0, n4570_o, n4563_o, n4556_o, n4549_o, n4542_o, n4535_o, n4528_o, n4521_o, n4514_o, n4507_o, n4500_o, n4493_o, n4486_o, n4479_o, n4472_o, n4465_o, n4451_o, n4458_o, n4444_o, 1'b0, 1'b0, n4435_o, n4425_o, n4415_o, n4405_o, n4395_o, n4385_o, n4375_o, n4365_o, n4355_o, n4345_o, n4335_o, n4325_o, n4315_o, n4305_o, n4295_o, n4285_o, mei_i, mti_i, msi_i};
  assign n4576_o = {21'b000000000000000000000, 21'b000000000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1500:16  */
  assign n4580_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1504:31  */
  assign n4583_o = trap_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1505:31  */
  assign n4585_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1506:31  */
  assign n4587_o = trap_ctrl[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1507:31  */
  assign n4589_o = trap_ctrl[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1507:108  */
  assign n4590_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1507:102  */
  assign n4592_o = {5'b00010, n4590_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1507:124  */
  assign n4593_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1507:118  */
  assign n4594_o = {n4592_o, n4593_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1508:31  */
  assign n4595_o = trap_ctrl[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1509:31  */
  assign n4597_o = trap_ctrl[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1510:31  */
  assign n4599_o = trap_ctrl[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1511:31  */
  assign n4601_o = trap_ctrl[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1512:31  */
  assign n4603_o = trap_ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1514:31  */
  assign n4605_o = trap_ctrl[52]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1515:31  */
  assign n4607_o = trap_ctrl[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1516:31  */
  assign n4609_o = trap_ctrl[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1517:31  */
  assign n4611_o = trap_ctrl[53]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1519:31  */
  assign n4613_o = trap_ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1520:31  */
  assign n4615_o = trap_ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1521:31  */
  assign n4617_o = trap_ctrl[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1522:31  */
  assign n4619_o = trap_ctrl[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1523:31  */
  assign n4621_o = trap_ctrl[40]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1524:31  */
  assign n4623_o = trap_ctrl[41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1525:31  */
  assign n4625_o = trap_ctrl[42]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1526:31  */
  assign n4627_o = trap_ctrl[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1527:31  */
  assign n4629_o = trap_ctrl[44]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1528:31  */
  assign n4631_o = trap_ctrl[45]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1529:31  */
  assign n4633_o = trap_ctrl[46]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1530:31  */
  assign n4635_o = trap_ctrl[47]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1531:31  */
  assign n4637_o = trap_ctrl[48]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1532:31  */
  assign n4639_o = trap_ctrl[49]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1533:31  */
  assign n4641_o = trap_ctrl[50]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1534:31  */
  assign n4643_o = trap_ctrl[51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1536:31  */
  assign n4645_o = trap_ctrl[35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1537:31  */
  assign n4647_o = trap_ctrl[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1537:7  */
  assign n4651_o = n4647_o ? 7'b1000011 : 7'b1000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1536:7  */
  assign n4652_o = n4645_o ? 7'b1001011 : n4651_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1534:7  */
  assign n4653_o = n4643_o ? 7'b1011111 : n4652_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1533:7  */
  assign n4654_o = n4641_o ? 7'b1011110 : n4653_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1532:7  */
  assign n4655_o = n4639_o ? 7'b1011101 : n4654_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1531:7  */
  assign n4656_o = n4637_o ? 7'b1011100 : n4655_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1530:7  */
  assign n4657_o = n4635_o ? 7'b1011011 : n4656_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1529:7  */
  assign n4658_o = n4633_o ? 7'b1011010 : n4657_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1528:7  */
  assign n4659_o = n4631_o ? 7'b1011001 : n4658_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1527:7  */
  assign n4660_o = n4629_o ? 7'b1011000 : n4659_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1526:7  */
  assign n4661_o = n4627_o ? 7'b1010111 : n4660_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1525:7  */
  assign n4662_o = n4625_o ? 7'b1010110 : n4661_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1524:7  */
  assign n4663_o = n4623_o ? 7'b1010101 : n4662_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1523:7  */
  assign n4664_o = n4621_o ? 7'b1010100 : n4663_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1522:7  */
  assign n4665_o = n4619_o ? 7'b1010011 : n4664_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1521:7  */
  assign n4666_o = n4617_o ? 7'b1010010 : n4665_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1520:7  */
  assign n4667_o = n4615_o ? 7'b1010001 : n4666_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1519:7  */
  assign n4668_o = n4613_o ? 7'b1010000 : n4667_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1517:7  */
  assign n4669_o = n4611_o ? 7'b1100100 : n4668_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1516:7  */
  assign n4670_o = n4609_o ? 7'b0100001 : n4669_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1515:7  */
  assign n4671_o = n4607_o ? 7'b0100010 : n4670_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1514:7  */
  assign n4672_o = n4605_o ? 7'b1100011 : n4671_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1512:7  */
  assign n4673_o = n4603_o ? 7'b0000101 : n4672_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1511:7  */
  assign n4674_o = n4601_o ? 7'b0000111 : n4673_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1510:7  */
  assign n4675_o = n4599_o ? 7'b0000100 : n4674_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1509:7  */
  assign n4676_o = n4597_o ? 7'b0000110 : n4675_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1508:7  */
  assign n4677_o = n4595_o ? 7'b0000011 : n4676_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1507:7  */
  assign n4678_o = n4589_o ? n4594_o : n4677_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1506:7  */
  assign n4679_o = n4587_o ? 7'b0000000 : n4678_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1505:7  */
  assign n4680_o = n4585_o ? 7'b0000010 : n4679_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1504:7  */
  assign n4681_o = n4583_o ? 7'b0000001 : n4680_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1549:16  */
  assign n4687_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1552:21  */
  assign n4690_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1552:33  */
  assign n4691_o = ~n4690_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1554:23  */
  assign n4692_o = trap_ctrl[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1554:54  */
  assign n4693_o = trap_ctrl[54]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1554:90  */
  assign n4694_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1554:96  */
  assign n4696_o = n4694_o == 4'b0110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1554:70  */
  assign n4697_o = n4696_o & n4693_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1554:39  */
  assign n4698_o = n4692_o | n4697_o;
  assign n4700_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1554:9  */
  assign n4701_o = n4698_o ? 1'b1 : n4700_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1557:24  */
  assign n4702_o = trap_ctrl[95]; // extract
  assign n4704_o = trap_ctrl[94]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1557:7  */
  assign n4705_o = n4702_o ? 1'b0 : n4704_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1552:7  */
  assign n4706_o = n4691_o ? n4701_o : n4705_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4718_o = trap_ctrl[53]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4720_o = 1'b0 | n4718_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4722_o = trap_ctrl[52]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4723_o = n4720_o | n4722_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4724_o = trap_ctrl[51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4725_o = n4723_o | n4724_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4726_o = trap_ctrl[50]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4727_o = n4725_o | n4726_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4728_o = trap_ctrl[49]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4729_o = n4727_o | n4728_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4730_o = trap_ctrl[48]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4731_o = n4729_o | n4730_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4732_o = trap_ctrl[47]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4733_o = n4731_o | n4732_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4734_o = trap_ctrl[46]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4735_o = n4733_o | n4734_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4736_o = trap_ctrl[45]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4737_o = n4735_o | n4736_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4738_o = trap_ctrl[44]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4739_o = n4737_o | n4738_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4740_o = trap_ctrl[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4741_o = n4739_o | n4740_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4742_o = trap_ctrl[42]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4743_o = n4741_o | n4742_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4744_o = trap_ctrl[41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4745_o = n4743_o | n4744_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4746_o = trap_ctrl[40]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4747_o = n4745_o | n4746_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4748_o = trap_ctrl[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4749_o = n4747_o | n4748_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4750_o = trap_ctrl[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4751_o = n4749_o | n4750_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4752_o = trap_ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4753_o = n4751_o | n4752_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4754_o = trap_ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4755_o = n4753_o | n4754_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4756_o = trap_ctrl[35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4757_o = n4755_o | n4756_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4758_o = trap_ctrl[34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4759_o = n4757_o | n4758_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4760_o = trap_ctrl[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4761_o = n4759_o | n4760_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1564:68  */
  assign n4762_o = debug_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1564:54  */
  assign n4763_o = n4761_o | n4762_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1564:83  */
  assign n4764_o = csr[339]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1564:76  */
  assign n4765_o = n4763_o | n4764_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4774_o = trap_ctrl[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4776_o = 1'b0 | n4774_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4778_o = trap_ctrl[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4779_o = n4776_o | n4778_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4780_o = trap_ctrl[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4781_o = n4779_o | n4780_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4782_o = trap_ctrl[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4783_o = n4781_o | n4782_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4784_o = trap_ctrl[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4785_o = n4783_o | n4784_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4786_o = trap_ctrl[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4787_o = n4785_o | n4786_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4788_o = trap_ctrl[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4789_o = n4787_o | n4788_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4790_o = trap_ctrl[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4791_o = n4789_o | n4790_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4792_o = trap_ctrl[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4793_o = n4791_o | n4792_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4794_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4795_o = n4793_o | n4794_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4796_o = trap_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4797_o = n4795_o | n4796_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1567:29  */
  assign n4798_o = n4797_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4808_o = trap_ctrl[51]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4810_o = 1'b0 | n4808_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4812_o = trap_ctrl[50]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4813_o = n4810_o | n4812_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4814_o = trap_ctrl[49]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4815_o = n4813_o | n4814_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4816_o = trap_ctrl[48]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4817_o = n4815_o | n4816_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4818_o = trap_ctrl[47]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4819_o = n4817_o | n4818_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4820_o = trap_ctrl[46]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4821_o = n4819_o | n4820_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4822_o = trap_ctrl[45]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4823_o = n4821_o | n4822_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4824_o = trap_ctrl[44]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4825_o = n4823_o | n4824_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4826_o = trap_ctrl[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4827_o = n4825_o | n4826_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4828_o = trap_ctrl[42]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4829_o = n4827_o | n4828_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4830_o = trap_ctrl[41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4831_o = n4829_o | n4830_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4832_o = trap_ctrl[40]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4833_o = n4831_o | n4832_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4834_o = trap_ctrl[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4835_o = n4833_o | n4834_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4836_o = trap_ctrl[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4837_o = n4835_o | n4836_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4838_o = trap_ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4839_o = n4837_o | n4838_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4840_o = trap_ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4841_o = n4839_o | n4840_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4842_o = trap_ctrl[35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4843_o = n4841_o | n4842_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4844_o = trap_ctrl[34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4845_o = n4843_o | n4844_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n4846_o = trap_ctrl[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n4847_o = n4845_o | n4846_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1573:12  */
  assign n4848_o = csr[127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1573:39  */
  assign n4849_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1573:49  */
  assign n4850_o = ~n4849_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1573:31  */
  assign n4851_o = n4848_o | n4850_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1572:81  */
  assign n4852_o = n4851_o & n4847_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1574:18  */
  assign n4853_o = debug_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1574:26  */
  assign n4854_o = ~n4853_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1573:67  */
  assign n4855_o = n4854_o & n4852_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1574:42  */
  assign n4856_o = csr[339]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1574:52  */
  assign n4857_o = ~n4856_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1574:33  */
  assign n4858_o = n4857_o & n4855_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1576:23  */
  assign n4859_o = trap_ctrl[53]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1575:7  */
  assign n4860_o = n4858_o | n4859_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1577:23  */
  assign n4861_o = trap_ctrl[52]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1576:46  */
  assign n4862_o = n4860_o | n4861_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1570:29  */
  assign n4863_o = n4862_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1580:35  */
  assign n4865_o = execute_engine[139:108]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1580:64  */
  assign n4866_o = trap_ctrl[61]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1580:43  */
  assign n4867_o = n4866_o ? n4865_o : n4868_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1580:114  */
  assign n4868_o = execute_engine[106:75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1589:33  */
  assign n4869_o = execute_engine[39:28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1591:24  */
  assign n4870_o = csr[11:10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1591:49  */
  assign n4871_o = csr[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1591:39  */
  assign n4872_o = {n4870_o, n4871_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1591:63  */
  assign n4873_o = csr[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1591:53  */
  assign n4874_o = {n4872_o, n4873_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1591:77  */
  assign n4875_o = csr[7:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1591:67  */
  assign n4876_o = {n4874_o, n4875_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1596:31  */
  assign n4877_o = execute_engine[22:20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1603:16  */
  assign n4880_o = csr[26]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1605:45  */
  assign n4881_o = execute_engine[27:23]; // extract
  assign n4883_o = n4882_o[31:5]; // extract
  assign n4884_o = {n4883_o, n4881_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1603:5  */
  assign n4885_o = n4880_o ? n4884_o : rs1_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1610:16  */
  assign n4886_o = csr[25:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1610:29  */
  assign n4888_o = n4886_o == 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1611:20  */
  assign n4889_o = ~n4885_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1610:5  */
  assign n4890_o = n4888_o ? n4889_o : n4885_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1618:15  */
  assign n4892_o = csr[25:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1619:9  */
  assign n4893_o = csr[94:63]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1619:23  */
  assign n4894_o = csr[126:95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1619:15  */
  assign n4895_o = n4893_o | n4894_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1619:29  */
  assign n4897_o = n4892_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1620:9  */
  assign n4898_o = csr[94:63]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1620:23  */
  assign n4899_o = csr[126:95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1620:15  */
  assign n4900_o = n4898_o & n4899_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1620:29  */
  assign n4902_o = n4892_o == 2'b11;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1621:23  */
  assign n4903_o = csr[126:95]; // extract
  assign n4904_o = {n4902_o, n4897_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1618:3  */
  always @*
    case (n4904_o)
      2'b10: n4905_o = n4900_o;
      2'b01: n4905_o = n4895_o;
      default: n4905_o = n4903_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1626:23  */
  assign n4906_o = csr[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1627:23  */
  assign n4907_o = csr[11:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1628:23  */
  assign n4908_o = csr[62:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1636:16  */
  assign n4910_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1670:21  */
  assign n4942_o = csr[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1670:54  */
  assign n4943_o = trap_ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1670:33  */
  assign n4944_o = ~n4943_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1670:28  */
  assign n4945_o = n4942_o & n4944_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:15  */
  assign n4946_o = csr[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:18  */
  assign n4947_o = csr[11:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1682:42  */
  assign n4948_o = csr[34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1683:42  */
  assign n4949_o = csr[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1685:44  */
  assign n4950_o = csr[42]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1685:61  */
  assign n4951_o = csr[43]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1685:49  */
  assign n4952_o = n4950_o | n4951_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1686:44  */
  assign n4953_o = csr[48]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1687:44  */
  assign n4954_o = csr[52]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1681:11  */
  assign n4956_o = n4947_o == 12'b001100000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1691:38  */
  assign n4957_o = csr[34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1692:38  */
  assign n4958_o = csr[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1693:38  */
  assign n4959_o = csr[42]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1694:38  */
  assign n4960_o = csr[62:47]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1690:11  */
  assign n4962_o = n4947_o == 12'b001100000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1697:26  */
  assign n4963_o = csr[32:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1697:39  */
  assign n4965_o = n4963_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1698:37  */
  assign n4966_o = csr[62:38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1698:55  */
  assign n4968_o = {n4966_o, 5'b00000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1698:65  */
  assign n4970_o = {n4968_o, 2'b01};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1700:37  */
  assign n4971_o = csr[62:33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1700:55  */
  assign n4973_o = {n4971_o, 2'b00};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1697:13  */
  assign n4974_o = n4965_o ? n4970_o : n4973_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1696:11  */
  assign n4976_o = n4947_o == 12'b001100000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1708:44  */
  assign n4977_o = csr[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1708:60  */
  assign n4978_o = csr[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1708:48  */
  assign n4979_o = n4977_o | n4978_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1703:11  */
  assign n4981_o = n4947_o == 12'b001100000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1718:33  */
  assign n4982_o = csr[62:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1717:11  */
  assign n4984_o = n4947_o == 12'b001101000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1721:34  */
  assign n4985_o = csr[62:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1721:52  */
  assign n4987_o = {n4985_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1720:11  */
  assign n4989_o = n4947_o == 12'b001101000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1727:36  */
  assign n4990_o = csr[62]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1727:52  */
  assign n4991_o = csr[35:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1727:41  */
  assign n4992_o = {n4990_o, n4991_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1726:11  */
  assign n4994_o = n4947_o == 12'b001101000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1737:48  */
  assign n4995_o = csr[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1738:48  */
  assign n4996_o = csr[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1735:11  */
  assign n4998_o = n4947_o == 12'b001100100000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1747:11  */
  assign n5000_o = n4947_o == 12'b011110110000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1757:11  */
  assign n5002_o = n4947_o == 12'b011110110001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1765:11  */
  assign n5004_o = n4947_o == 12'b011110110010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1773:11  */
  assign n5006_o = n4947_o == 12'b011110100001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1784:11  */
  assign n5008_o = n4947_o == 12'b011110100010;
  assign n5009_o = {n5008_o, n5006_o, n5004_o, n5002_o, n5000_o, n4998_o, n4994_o, n4989_o, n4984_o, n4981_o, n4976_o, n4962_o, n4956_o};
  assign n5010_o = csr[127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5011_o = n5010_o;
      13'b0100000000000: n5011_o = n5010_o;
      13'b0010000000000: n5011_o = n5010_o;
      13'b0001000000000: n5011_o = n5010_o;
      13'b0000100000000: n5011_o = n5010_o;
      13'b0000010000000: n5011_o = n5010_o;
      13'b0000001000000: n5011_o = n5010_o;
      13'b0000000100000: n5011_o = n5010_o;
      13'b0000000010000: n5011_o = n5010_o;
      13'b0000000001000: n5011_o = n5010_o;
      13'b0000000000100: n5011_o = n5010_o;
      13'b0000000000010: n5011_o = n5010_o;
      13'b0000000000001: n5011_o = n4948_o;
      default: n5011_o = n5010_o;
    endcase
  assign n5012_o = csr[128]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5013_o = n5012_o;
      13'b0100000000000: n5013_o = n5012_o;
      13'b0010000000000: n5013_o = n5012_o;
      13'b0001000000000: n5013_o = n5012_o;
      13'b0000100000000: n5013_o = n5012_o;
      13'b0000010000000: n5013_o = n5012_o;
      13'b0000001000000: n5013_o = n5012_o;
      13'b0000000100000: n5013_o = n5012_o;
      13'b0000000010000: n5013_o = n5012_o;
      13'b0000000001000: n5013_o = n5012_o;
      13'b0000000000100: n5013_o = n5012_o;
      13'b0000000000010: n5013_o = n5012_o;
      13'b0000000000001: n5013_o = n4949_o;
      default: n5013_o = n5012_o;
    endcase
  assign n5014_o = csr[129]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5015_o = n5014_o;
      13'b0100000000000: n5015_o = n5014_o;
      13'b0010000000000: n5015_o = n5014_o;
      13'b0001000000000: n5015_o = n5014_o;
      13'b0000100000000: n5015_o = n5014_o;
      13'b0000010000000: n5015_o = n5014_o;
      13'b0000001000000: n5015_o = n5014_o;
      13'b0000000100000: n5015_o = n5014_o;
      13'b0000000010000: n5015_o = n5014_o;
      13'b0000000001000: n5015_o = n5014_o;
      13'b0000000000100: n5015_o = n5014_o;
      13'b0000000000010: n5015_o = n5014_o;
      13'b0000000000001: n5015_o = n4952_o;
      default: n5015_o = n5014_o;
    endcase
  assign n5016_o = csr[130]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5017_o = n5016_o;
      13'b0100000000000: n5017_o = n5016_o;
      13'b0010000000000: n5017_o = n5016_o;
      13'b0001000000000: n5017_o = n5016_o;
      13'b0000100000000: n5017_o = n5016_o;
      13'b0000010000000: n5017_o = n5016_o;
      13'b0000001000000: n5017_o = n5016_o;
      13'b0000000100000: n5017_o = n5016_o;
      13'b0000000010000: n5017_o = n5016_o;
      13'b0000000001000: n5017_o = n5016_o;
      13'b0000000000100: n5017_o = n5016_o;
      13'b0000000000010: n5017_o = n5016_o;
      13'b0000000000001: n5017_o = n4953_o;
      default: n5017_o = n5016_o;
    endcase
  assign n5018_o = csr[131]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5019_o = n5018_o;
      13'b0100000000000: n5019_o = n5018_o;
      13'b0010000000000: n5019_o = n5018_o;
      13'b0001000000000: n5019_o = n5018_o;
      13'b0000100000000: n5019_o = n5018_o;
      13'b0000010000000: n5019_o = n5018_o;
      13'b0000001000000: n5019_o = n5018_o;
      13'b0000000100000: n5019_o = n5018_o;
      13'b0000000010000: n5019_o = n5018_o;
      13'b0000000001000: n5019_o = n5018_o;
      13'b0000000000100: n5019_o = n5018_o;
      13'b0000000000010: n5019_o = n5018_o;
      13'b0000000000001: n5019_o = n4954_o;
      default: n5019_o = n5018_o;
    endcase
  assign n5020_o = csr[132]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5021_o = n5020_o;
      13'b0100000000000: n5021_o = n5020_o;
      13'b0010000000000: n5021_o = n5020_o;
      13'b0001000000000: n5021_o = n5020_o;
      13'b0000100000000: n5021_o = n5020_o;
      13'b0000010000000: n5021_o = n5020_o;
      13'b0000001000000: n5021_o = n5020_o;
      13'b0000000100000: n5021_o = n5020_o;
      13'b0000000010000: n5021_o = n5020_o;
      13'b0000000001000: n5021_o = n5020_o;
      13'b0000000000100: n5021_o = n5020_o;
      13'b0000000000010: n5021_o = n4957_o;
      13'b0000000000001: n5021_o = n5020_o;
      default: n5021_o = n5020_o;
    endcase
  assign n5022_o = csr[133]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5023_o = n5022_o;
      13'b0100000000000: n5023_o = n5022_o;
      13'b0010000000000: n5023_o = n5022_o;
      13'b0001000000000: n5023_o = n5022_o;
      13'b0000100000000: n5023_o = n5022_o;
      13'b0000010000000: n5023_o = n5022_o;
      13'b0000001000000: n5023_o = n5022_o;
      13'b0000000100000: n5023_o = n5022_o;
      13'b0000000010000: n5023_o = n5022_o;
      13'b0000000001000: n5023_o = n5022_o;
      13'b0000000000100: n5023_o = n5022_o;
      13'b0000000000010: n5023_o = n4959_o;
      13'b0000000000001: n5023_o = n5022_o;
      default: n5023_o = n5022_o;
    endcase
  assign n5024_o = csr[134]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5025_o = n5024_o;
      13'b0100000000000: n5025_o = n5024_o;
      13'b0010000000000: n5025_o = n5024_o;
      13'b0001000000000: n5025_o = n5024_o;
      13'b0000100000000: n5025_o = n5024_o;
      13'b0000010000000: n5025_o = n5024_o;
      13'b0000001000000: n5025_o = n5024_o;
      13'b0000000100000: n5025_o = n5024_o;
      13'b0000000010000: n5025_o = n5024_o;
      13'b0000000001000: n5025_o = n5024_o;
      13'b0000000000100: n5025_o = n5024_o;
      13'b0000000000010: n5025_o = n4958_o;
      13'b0000000000001: n5025_o = n5024_o;
      default: n5025_o = n5024_o;
    endcase
  assign n5026_o = csr[150:135]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5027_o = n5026_o;
      13'b0100000000000: n5027_o = n5026_o;
      13'b0010000000000: n5027_o = n5026_o;
      13'b0001000000000: n5027_o = n5026_o;
      13'b0000100000000: n5027_o = n5026_o;
      13'b0000010000000: n5027_o = n5026_o;
      13'b0000001000000: n5027_o = n5026_o;
      13'b0000000100000: n5027_o = n5026_o;
      13'b0000000010000: n5027_o = n5026_o;
      13'b0000000001000: n5027_o = n5026_o;
      13'b0000000000100: n5027_o = n5026_o;
      13'b0000000000010: n5027_o = n4960_o;
      13'b0000000000001: n5027_o = n5026_o;
      default: n5027_o = n5026_o;
    endcase
  assign n5028_o = csr[185:154]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5029_o = n5028_o;
      13'b0100000000000: n5029_o = n5028_o;
      13'b0010000000000: n5029_o = n5028_o;
      13'b0001000000000: n5029_o = n5028_o;
      13'b0000100000000: n5029_o = n5028_o;
      13'b0000010000000: n5029_o = n5028_o;
      13'b0000001000000: n5029_o = n5028_o;
      13'b0000000100000: n5029_o = n4987_o;
      13'b0000000010000: n5029_o = n5028_o;
      13'b0000000001000: n5029_o = n5028_o;
      13'b0000000000100: n5029_o = n5028_o;
      13'b0000000000010: n5029_o = n5028_o;
      13'b0000000000001: n5029_o = n5028_o;
      default: n5029_o = n5028_o;
    endcase
  assign n5030_o = csr[191:186]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5031_o = n5030_o;
      13'b0100000000000: n5031_o = n5030_o;
      13'b0010000000000: n5031_o = n5030_o;
      13'b0001000000000: n5031_o = n5030_o;
      13'b0000100000000: n5031_o = n5030_o;
      13'b0000010000000: n5031_o = n5030_o;
      13'b0000001000000: n5031_o = n4992_o;
      13'b0000000100000: n5031_o = n5030_o;
      13'b0000000010000: n5031_o = n5030_o;
      13'b0000000001000: n5031_o = n5030_o;
      13'b0000000000100: n5031_o = n5030_o;
      13'b0000000000010: n5031_o = n5030_o;
      13'b0000000000001: n5031_o = n5030_o;
      default: n5031_o = n5030_o;
    endcase
  assign n5032_o = csr[223:192]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5033_o = n5032_o;
      13'b0100000000000: n5033_o = n5032_o;
      13'b0010000000000: n5033_o = n5032_o;
      13'b0001000000000: n5033_o = n5032_o;
      13'b0000100000000: n5033_o = n5032_o;
      13'b0000010000000: n5033_o = n5032_o;
      13'b0000001000000: n5033_o = n5032_o;
      13'b0000000100000: n5033_o = n5032_o;
      13'b0000000010000: n5033_o = n5032_o;
      13'b0000000001000: n5033_o = n5032_o;
      13'b0000000000100: n5033_o = n4974_o;
      13'b0000000000010: n5033_o = n5032_o;
      13'b0000000000001: n5033_o = n5032_o;
      default: n5033_o = n5032_o;
    endcase
  assign n5034_o = csr[319:288]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5035_o = n5034_o;
      13'b0100000000000: n5035_o = n5034_o;
      13'b0010000000000: n5035_o = n5034_o;
      13'b0001000000000: n5035_o = n5034_o;
      13'b0000100000000: n5035_o = n5034_o;
      13'b0000010000000: n5035_o = n5034_o;
      13'b0000001000000: n5035_o = n5034_o;
      13'b0000000100000: n5035_o = n5034_o;
      13'b0000000010000: n5035_o = n4982_o;
      13'b0000000001000: n5035_o = n5034_o;
      13'b0000000000100: n5035_o = n5034_o;
      13'b0000000000010: n5035_o = n5034_o;
      13'b0000000000001: n5035_o = n5034_o;
      default: n5035_o = n5034_o;
    endcase
  assign n5036_o = csr[320]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5037_o = n5036_o;
      13'b0100000000000: n5037_o = n5036_o;
      13'b0010000000000: n5037_o = n5036_o;
      13'b0001000000000: n5037_o = n5036_o;
      13'b0000100000000: n5037_o = n5036_o;
      13'b0000010000000: n5037_o = n5036_o;
      13'b0000001000000: n5037_o = n5036_o;
      13'b0000000100000: n5037_o = n5036_o;
      13'b0000000010000: n5037_o = n5036_o;
      13'b0000000001000: n5037_o = n4979_o;
      13'b0000000000100: n5037_o = n5036_o;
      13'b0000000000010: n5037_o = n5036_o;
      13'b0000000000001: n5037_o = n5036_o;
      default: n5037_o = n5036_o;
    endcase
  assign n5038_o = csr[321]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5039_o = n5038_o;
      13'b0100000000000: n5039_o = n5038_o;
      13'b0010000000000: n5039_o = n5038_o;
      13'b0001000000000: n5039_o = n5038_o;
      13'b0000100000000: n5039_o = n5038_o;
      13'b0000010000000: n5039_o = n4995_o;
      13'b0000001000000: n5039_o = n5038_o;
      13'b0000000100000: n5039_o = n5038_o;
      13'b0000000010000: n5039_o = n5038_o;
      13'b0000000001000: n5039_o = n5038_o;
      13'b0000000000100: n5039_o = n5038_o;
      13'b0000000000010: n5039_o = n5038_o;
      13'b0000000000001: n5039_o = n5038_o;
      default: n5039_o = n5038_o;
    endcase
  assign n5040_o = csr[323]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1676:9  */
  always @*
    case (n5009_o)
      13'b1000000000000: n5041_o = n5040_o;
      13'b0100000000000: n5041_o = n5040_o;
      13'b0010000000000: n5041_o = n5040_o;
      13'b0001000000000: n5041_o = n5040_o;
      13'b0000100000000: n5041_o = n5040_o;
      13'b0000010000000: n5041_o = n4996_o;
      13'b0000001000000: n5041_o = n5040_o;
      13'b0000000100000: n5041_o = n5040_o;
      13'b0000000010000: n5041_o = n5040_o;
      13'b0000000001000: n5041_o = n5040_o;
      13'b0000000000100: n5041_o = n5040_o;
      13'b0000000000010: n5041_o = n5040_o;
      13'b0000000000001: n5041_o = n5040_o;
      default: n5041_o = n5040_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1801:24  */
  assign n5042_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1805:40  */
  assign n5043_o = trap_ctrl[61]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1805:80  */
  assign n5044_o = trap_ctrl[59:55]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1805:63  */
  assign n5045_o = {n5043_o, n5044_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1806:38  */
  assign n5046_o = trap_ctrl[93:63]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1806:56  */
  assign n5048_o = {n5046_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1808:30  */
  assign n5049_o = trap_ctrl[61]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1808:34  */
  assign n5050_o = ~n5049_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1808:61  */
  assign n5051_o = trap_ctrl[57]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1808:41  */
  assign n5052_o = n5051_o & n5050_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1808:11  */
  assign n5054_o = n5052_o ? mar_i : 32'b00000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1814:30  */
  assign n5055_o = trap_ctrl[61]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1814:34  */
  assign n5056_o = ~n5055_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1816:32  */
  assign n5058_o = execute_engine[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1816:45  */
  assign n5060_o = 1'b1 & n5058_o;
  assign n5062_o = execute_engine[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1816:13  */
  assign n5063_o = n5060_o ? 1'b0 : n5062_o;
  assign n5064_o = execute_engine[39:10]; // extract
  assign n5065_o = execute_engine[8]; // extract
  assign n5067_o = {n5064_o, n5063_o, n5065_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1814:11  */
  assign n5068_o = n5056_o ? n5067_o : 32'b00000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1825:35  */
  assign n5071_o = csr[127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1826:35  */
  assign n5072_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1842:24  */
  assign n5073_o = trap_ctrl[96]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1856:36  */
  assign n5074_o = csr[129]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1858:21  */
  assign n5076_o = csr[129]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1858:33  */
  assign n5078_o = n5076_o != 1'b1;
  assign n5080_o = csr[130]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1858:13  */
  assign n5081_o = n5078_o ? 1'b0 : n5080_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1862:35  */
  assign n5082_o = csr[128]; // extract
  assign n5084_o = {n5081_o, 1'b0, 1'b1, n5082_o};
  assign n5085_o = csr[130:127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1842:7  */
  assign n5086_o = n5073_o ? n5084_o : n5085_o;
  assign n5087_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1842:7  */
  assign n5088_o = n5073_o ? n5074_o : n5087_o;
  assign n5089_o = {n5072_o, n5071_o, 1'b0};
  assign n5090_o = {n5045_o, n5048_o};
  assign n5091_o = {n5068_o, n5054_o};
  assign n5092_o = n5086_o[2:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1801:7  */
  assign n5093_o = n5042_o ? n5089_o : n5092_o;
  assign n5094_o = n5086_o[3]; // extract
  assign n5095_o = csr[130]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1801:7  */
  assign n5096_o = n5042_o ? n5095_o : n5094_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1801:7  */
  assign n5097_o = n5042_o ? 1'b1 : n5088_o;
  assign n5098_o = csr[191:154]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1801:7  */
  assign n5099_o = n5042_o ? n5090_o : n5098_o;
  assign n5100_o = csr[287:224]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1801:7  */
  assign n5101_o = n5042_o ? n5091_o : n5100_o;
  assign n5102_o = {n5096_o, n5093_o};
  assign n5103_o = {n5027_o, n5025_o, n5023_o, n5021_o, n5019_o, n5017_o, n5015_o, n5013_o, n5011_o};
  assign n5104_o = {n5033_o, n5031_o, n5029_o};
  assign n5105_o = {n5039_o, n5037_o, n5035_o};
  assign n5106_o = n5103_o[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:7  */
  assign n5107_o = n4946_o ? n5106_o : n5102_o;
  assign n5108_o = n5103_o[23:4]; // extract
  assign n5109_o = csr[150:131]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:7  */
  assign n5110_o = n4946_o ? n5108_o : n5109_o;
  assign n5111_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:7  */
  assign n5112_o = n4946_o ? n5111_o : n5097_o;
  assign n5113_o = n5104_o[37:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:7  */
  assign n5114_o = n4946_o ? n5113_o : n5099_o;
  assign n5115_o = n5104_o[69:38]; // extract
  assign n5116_o = csr[223:192]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:7  */
  assign n5117_o = n4946_o ? n5115_o : n5116_o;
  assign n5118_o = csr[287:224]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:7  */
  assign n5119_o = n4946_o ? n5118_o : n5101_o;
  assign n5120_o = csr[321:288]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:7  */
  assign n5121_o = n4946_o ? n5105_o : n5120_o;
  assign n5122_o = csr[323]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1675:7  */
  assign n5123_o = n4946_o ? n5041_o : n5122_o;
  assign n5137_o = {n5110_o, n5107_o};
  assign n5138_o = {3'b000, 1'b1, 1'b0, 1'b0, 1'b0, 13'b0000000000000, n5123_o, 1'b0, n5121_o, n5119_o, n5117_o, n5114_o};
  assign n5139_o = {32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  assign n5140_o = {1'b0, 1'b0, 1'b0};
  assign n5155_o = {16'b0000000000000000, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
  assign n5156_o = {3'b000, 1'b1, 1'b0, 1'b0, 1'b0, 16'b0000000000000000, 1'b0, 32'b00011001100010000000011100000100, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 6'b000000, 32'b00000000000000000000000000000000};
  assign n5157_o = {32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  assign n5158_o = {1'b0, 1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1924:38  */
  assign n5168_o = csr[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1924:60  */
  assign n5169_o = csr[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1924:48  */
  assign n5170_o = n5169_o & n5168_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1924:80  */
  assign n5171_o = csr[11:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1924:85  */
  assign n5173_o = n5171_o == 12'b001101000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1924:71  */
  assign n5174_o = n5173_o & n5170_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1924:28  */
  assign n5175_o = n5174_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1925:38  */
  assign n5178_o = csr[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1925:60  */
  assign n5179_o = csr[24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1925:48  */
  assign n5180_o = n5179_o & n5178_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1925:80  */
  assign n5181_o = csr[11:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1925:85  */
  assign n5183_o = n5181_o == 12'b011110100001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1925:71  */
  assign n5184_o = n5183_o & n5180_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1925:28  */
  assign n5185_o = n5184_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1928:55  */
  assign n5188_o = debug_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1928:38  */
  assign n5189_o = n5188_o ? 1'b1 : n5190_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1928:79  */
  assign n5190_o = csr[152]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:14  */
  assign n5192_o = csr[23:12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1942:30  */
  assign n5193_o = csr[127]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1943:30  */
  assign n5194_o = csr[128]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1944:51  */
  assign n5195_o = csr[129]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1944:51  */
  assign n5196_o = csr[129]; // extract
  assign n5197_o = {n5195_o, n5196_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1945:30  */
  assign n5198_o = csr[130]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1946:30  */
  assign n5199_o = csr[131]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1946:41  */
  assign n5202_o = n5199_o & 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1941:7  */
  assign n5204_o = n5192_o == 12'b001100000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1950:7  */
  assign n5222_o = n5192_o == 12'b001100000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1962:30  */
  assign n5223_o = csr[132]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1963:30  */
  assign n5224_o = csr[134]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1964:30  */
  assign n5225_o = csr[133]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1965:40  */
  assign n5226_o = csr[150:135]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1961:7  */
  assign n5228_o = n5192_o == 12'b001100000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1968:26  */
  assign n5229_o = csr[223:192]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1967:7  */
  assign n5231_o = n5192_o == 12'b001100000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1973:33  */
  assign n5232_o = csr[320]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1974:33  */
  assign n5233_o = csr[320]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1970:7  */
  assign n5235_o = n5192_o == 12'b001100000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1991:26  */
  assign n5236_o = csr[319:288]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1990:7  */
  assign n5238_o = n5192_o == 12'b001101000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1994:30  */
  assign n5239_o = csr[185:155]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1994:48  */
  assign n5241_o = {n5239_o, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1993:7  */
  assign n5243_o = n5192_o == 12'b001101000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1997:44  */
  assign n5244_o = csr[191]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1998:44  */
  assign n5245_o = csr[190:186]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1996:7  */
  assign n5247_o = n5192_o == 12'b001101000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2001:26  */
  assign n5248_o = csr[255:224]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2000:7  */
  assign n5250_o = n5192_o == 12'b001101000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2004:53  */
  assign n5251_o = trap_ctrl[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2005:53  */
  assign n5252_o = trap_ctrl[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2006:53  */
  assign n5253_o = trap_ctrl[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2007:53  */
  assign n5254_o = trap_ctrl[30:15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2003:7  */
  assign n5256_o = n5192_o == 12'b001101000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2010:26  */
  assign n5257_o = csr[287:256]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2009:7  */
  assign n5259_o = n5192_o == 12'b001101001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2017:44  */
  assign n5260_o = csr[321]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2018:44  */
  assign n5261_o = csr[323]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2015:7  */
  assign n5263_o = n5192_o == 12'b001100100000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2027:7  */
  assign n5265_o = n5192_o == 12'b001100100011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2028:7  */
  assign n5267_o = n5192_o == 12'b001100100100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2029:7  */
  assign n5269_o = n5192_o == 12'b001100100101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2030:7  */
  assign n5271_o = n5192_o == 12'b001100100110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2031:7  */
  assign n5273_o = n5192_o == 12'b001100100111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2032:7  */
  assign n5275_o = n5192_o == 12'b001100101000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2033:7  */
  assign n5277_o = n5192_o == 12'b001100101001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2034:7  */
  assign n5279_o = n5192_o == 12'b001100101010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2035:7  */
  assign n5281_o = n5192_o == 12'b001100101011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2036:7  */
  assign n5283_o = n5192_o == 12'b001100101100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2037:7  */
  assign n5285_o = n5192_o == 12'b001100101101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2038:7  */
  assign n5287_o = n5192_o == 12'b001100101110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2039:7  */
  assign n5289_o = n5192_o == 12'b001100101111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2045:115  */
  assign n5290_o = cnt_lo_rd[95:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2045:7  */
  assign n5292_o = n5192_o == 12'b101100000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2045:32  */
  assign n5294_o = n5192_o == 12'b110000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2045:32  */
  assign n5295_o = n5292_o | n5294_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2046:115  */
  assign n5296_o = cnt_lo_rd[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2046:7  */
  assign n5298_o = n5192_o == 12'b101100000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2046:32  */
  assign n5300_o = n5192_o == 12'b110000000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2046:32  */
  assign n5301_o = n5298_o | n5300_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2047:7  */
  assign n5303_o = n5192_o == 12'b101100000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2047:32  */
  assign n5305_o = n5192_o == 12'b110000000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2047:32  */
  assign n5306_o = n5303_o | n5305_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2048:7  */
  assign n5308_o = n5192_o == 12'b101100000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2048:32  */
  assign n5310_o = n5192_o == 12'b110000000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2048:32  */
  assign n5311_o = n5308_o | n5310_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2049:7  */
  assign n5313_o = n5192_o == 12'b101100000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2049:32  */
  assign n5315_o = n5192_o == 12'b110000000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2049:32  */
  assign n5316_o = n5313_o | n5315_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2050:7  */
  assign n5318_o = n5192_o == 12'b101100000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2050:32  */
  assign n5320_o = n5192_o == 12'b110000000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2050:32  */
  assign n5321_o = n5318_o | n5320_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2051:7  */
  assign n5323_o = n5192_o == 12'b101100000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2051:32  */
  assign n5325_o = n5192_o == 12'b110000000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2051:32  */
  assign n5326_o = n5323_o | n5325_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2052:7  */
  assign n5328_o = n5192_o == 12'b101100001000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2052:32  */
  assign n5330_o = n5192_o == 12'b110000001000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2052:32  */
  assign n5331_o = n5328_o | n5330_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2053:7  */
  assign n5333_o = n5192_o == 12'b101100001001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2053:32  */
  assign n5335_o = n5192_o == 12'b110000001001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2053:32  */
  assign n5336_o = n5333_o | n5335_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2054:7  */
  assign n5338_o = n5192_o == 12'b101100001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2054:32  */
  assign n5340_o = n5192_o == 12'b110000001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2054:32  */
  assign n5341_o = n5338_o | n5340_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2055:7  */
  assign n5343_o = n5192_o == 12'b101100001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2055:32  */
  assign n5345_o = n5192_o == 12'b110000001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2055:32  */
  assign n5346_o = n5343_o | n5345_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2056:7  */
  assign n5348_o = n5192_o == 12'b101100001100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2056:32  */
  assign n5350_o = n5192_o == 12'b110000001100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2056:32  */
  assign n5351_o = n5348_o | n5350_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2057:7  */
  assign n5353_o = n5192_o == 12'b101100001101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2057:32  */
  assign n5355_o = n5192_o == 12'b110000001101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2057:32  */
  assign n5356_o = n5353_o | n5355_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2058:7  */
  assign n5358_o = n5192_o == 12'b101100001110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2058:32  */
  assign n5360_o = n5192_o == 12'b110000001110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2058:32  */
  assign n5361_o = n5358_o | n5360_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2059:7  */
  assign n5363_o = n5192_o == 12'b101100001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2059:32  */
  assign n5365_o = n5192_o == 12'b110000001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2059:32  */
  assign n5366_o = n5363_o | n5365_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2062:117  */
  assign n5367_o = cnt_hi_rd[95:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2062:7  */
  assign n5369_o = n5192_o == 12'b101110000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2062:33  */
  assign n5371_o = n5192_o == 12'b110010000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2062:33  */
  assign n5372_o = n5369_o | n5371_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2063:117  */
  assign n5373_o = cnt_hi_rd[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2063:7  */
  assign n5375_o = n5192_o == 12'b101110000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2063:33  */
  assign n5377_o = n5192_o == 12'b110010000010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2063:33  */
  assign n5378_o = n5375_o | n5377_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2064:7  */
  assign n5380_o = n5192_o == 12'b101110000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2064:33  */
  assign n5382_o = n5192_o == 12'b110010000011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2064:33  */
  assign n5383_o = n5380_o | n5382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2065:7  */
  assign n5385_o = n5192_o == 12'b101110000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2065:33  */
  assign n5387_o = n5192_o == 12'b110010000100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2065:33  */
  assign n5388_o = n5385_o | n5387_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2066:7  */
  assign n5390_o = n5192_o == 12'b101110000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2066:33  */
  assign n5392_o = n5192_o == 12'b110010000101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2066:33  */
  assign n5393_o = n5390_o | n5392_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2067:7  */
  assign n5395_o = n5192_o == 12'b101110000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2067:33  */
  assign n5397_o = n5192_o == 12'b110010000110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2067:33  */
  assign n5398_o = n5395_o | n5397_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2068:7  */
  assign n5400_o = n5192_o == 12'b101110000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2068:33  */
  assign n5402_o = n5192_o == 12'b110010000111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2068:33  */
  assign n5403_o = n5400_o | n5402_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2069:7  */
  assign n5405_o = n5192_o == 12'b101110001000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2069:33  */
  assign n5407_o = n5192_o == 12'b110010001000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2069:33  */
  assign n5408_o = n5405_o | n5407_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2070:7  */
  assign n5410_o = n5192_o == 12'b101110001001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2070:33  */
  assign n5412_o = n5192_o == 12'b110010001001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2070:33  */
  assign n5413_o = n5410_o | n5412_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2071:7  */
  assign n5415_o = n5192_o == 12'b101110001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2071:33  */
  assign n5417_o = n5192_o == 12'b110010001010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2071:33  */
  assign n5418_o = n5415_o | n5417_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2072:7  */
  assign n5420_o = n5192_o == 12'b101110001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2072:33  */
  assign n5422_o = n5192_o == 12'b110010001011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2072:33  */
  assign n5423_o = n5420_o | n5422_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2073:7  */
  assign n5425_o = n5192_o == 12'b101110001100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2073:33  */
  assign n5427_o = n5192_o == 12'b110010001100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2073:33  */
  assign n5428_o = n5425_o | n5427_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2074:7  */
  assign n5430_o = n5192_o == 12'b101110001101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2074:33  */
  assign n5432_o = n5192_o == 12'b110010001101;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2074:33  */
  assign n5433_o = n5430_o | n5432_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2075:7  */
  assign n5435_o = n5192_o == 12'b101110001110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2075:33  */
  assign n5437_o = n5192_o == 12'b110010001110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2075:33  */
  assign n5438_o = n5435_o | n5437_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2076:7  */
  assign n5440_o = n5192_o == 12'b101110001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2076:33  */
  assign n5442_o = n5192_o == 12'b110010001111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2076:33  */
  assign n5443_o = n5440_o | n5442_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2081:7  */
  assign n5445_o = n5192_o == 12'b111100010001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2082:7  */
  assign n5448_o = n5192_o == 12'b111100010010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2083:7  */
  assign n5450_o = n5192_o == 12'b111100010011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2084:7  */
  assign n5452_o = n5192_o == 12'b111100010100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2090:7  */
  assign n5454_o = n5192_o == 12'b011110110000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2091:7  */
  assign n5456_o = n5192_o == 12'b011110110001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2092:7  */
  assign n5458_o = n5192_o == 12'b011110110010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2098:7  */
  assign n5460_o = n5192_o == 12'b011110100001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2099:7  */
  assign n5462_o = n5192_o == 12'b011110100010;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2100:7  */
  assign n5464_o = n5192_o == 12'b011110100100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2110:7  */
  assign n5495_o = n5192_o == 12'b111111000000;
  assign n5496_o = {n5495_o, n5464_o, n5462_o, n5460_o, n5458_o, n5456_o, n5454_o, n5452_o, n5450_o, n5448_o, n5445_o, n5443_o, n5438_o, n5433_o, n5428_o, n5423_o, n5418_o, n5413_o, n5408_o, n5403_o, n5398_o, n5393_o, n5388_o, n5383_o, n5378_o, n5372_o, n5366_o, n5361_o, n5356_o, n5351_o, n5346_o, n5341_o, n5336_o, n5331_o, n5326_o, n5321_o, n5316_o, n5311_o, n5306_o, n5301_o, n5295_o, n5289_o, n5287_o, n5285_o, n5283_o, n5281_o, n5279_o, n5277_o, n5275_o, n5273_o, n5271_o, n5269_o, n5267_o, n5265_o, n5263_o, n5259_o, n5256_o, n5250_o, n5247_o, n5243_o, n5238_o, n5235_o, n5231_o, n5228_o, n5222_o, n5204_o};
  assign n5497_o = n5229_o[0]; // extract
  assign n5498_o = n5236_o[0]; // extract
  assign n5499_o = n5241_o[0]; // extract
  assign n5500_o = n5245_o[0]; // extract
  assign n5501_o = n5248_o[0]; // extract
  assign n5502_o = n5257_o[0]; // extract
  assign n5503_o = n5290_o[0]; // extract
  assign n5504_o = n5296_o[0]; // extract
  assign n5505_o = n5367_o[0]; // extract
  assign n5506_o = n5373_o[0]; // extract
  assign n5508_o = n5446_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b1;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5512_o = n5508_o;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5512_o = n5506_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5512_o = n5505_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5512_o = n5504_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5512_o = n5503_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5512_o = n5260_o;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5512_o = n5502_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5512_o = n5501_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5512_o = n5500_o;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5512_o = n5499_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5512_o = n5498_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5512_o = n5232_o;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5512_o = n5497_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5512_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5512_o = 1'b0;
      default: n5512_o = 1'b0;
    endcase
  assign n5513_o = n5229_o[1]; // extract
  assign n5514_o = n5236_o[1]; // extract
  assign n5515_o = n5241_o[1]; // extract
  assign n5516_o = n5245_o[1]; // extract
  assign n5517_o = n5248_o[1]; // extract
  assign n5518_o = n5257_o[1]; // extract
  assign n5519_o = n5290_o[1]; // extract
  assign n5520_o = n5296_o[1]; // extract
  assign n5521_o = n5367_o[1]; // extract
  assign n5522_o = n5373_o[1]; // extract
  assign n5524_o = n5446_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b1;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5528_o = n5524_o;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5528_o = n5522_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5528_o = n5521_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5528_o = n5520_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5528_o = n5519_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5528_o = n5518_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5528_o = n5517_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5528_o = n5516_o;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5528_o = n5515_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5528_o = n5514_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5528_o = n5513_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5528_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5528_o = 1'b0;
      default: n5528_o = 1'b0;
    endcase
  assign n5529_o = n5229_o[2]; // extract
  assign n5530_o = n5236_o[2]; // extract
  assign n5531_o = n5241_o[2]; // extract
  assign n5532_o = n5245_o[2]; // extract
  assign n5533_o = n5248_o[2]; // extract
  assign n5534_o = n5257_o[2]; // extract
  assign n5535_o = n5290_o[2]; // extract
  assign n5536_o = n5296_o[2]; // extract
  assign n5537_o = n5367_o[2]; // extract
  assign n5538_o = n5373_o[2]; // extract
  assign n5540_o = n5446_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5544_o = n5540_o;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5544_o = n5538_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5544_o = n5537_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5544_o = n5536_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5544_o = n5535_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5544_o = n5261_o;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5544_o = n5534_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5544_o = n5533_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5544_o = n5532_o;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5544_o = n5531_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5544_o = n5530_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5544_o = n5233_o;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5544_o = n5529_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5544_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5544_o = 1'b1;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5544_o = 1'b0;
      default: n5544_o = 1'b0;
    endcase
  assign n5545_o = n5229_o[3]; // extract
  assign n5546_o = n5236_o[3]; // extract
  assign n5547_o = n5241_o[3]; // extract
  assign n5548_o = n5245_o[3]; // extract
  assign n5549_o = n5248_o[3]; // extract
  assign n5550_o = n5257_o[3]; // extract
  assign n5551_o = n5290_o[3]; // extract
  assign n5552_o = n5296_o[3]; // extract
  assign n5553_o = n5367_o[3]; // extract
  assign n5554_o = n5373_o[3]; // extract
  assign n5556_o = n5446_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5560_o = n5556_o;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5560_o = n5554_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5560_o = n5553_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5560_o = n5552_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5560_o = n5551_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5560_o = n5550_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5560_o = n5251_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5560_o = n5549_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5560_o = n5548_o;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5560_o = n5547_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5560_o = n5546_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5560_o = n5545_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5560_o = n5223_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5560_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5560_o = n5193_o;
      default: n5560_o = 1'b0;
    endcase
  assign n5561_o = n5229_o[4]; // extract
  assign n5562_o = n5236_o[4]; // extract
  assign n5563_o = n5241_o[4]; // extract
  assign n5564_o = n5245_o[4]; // extract
  assign n5565_o = n5248_o[4]; // extract
  assign n5566_o = n5257_o[4]; // extract
  assign n5567_o = n5290_o[4]; // extract
  assign n5568_o = n5296_o[4]; // extract
  assign n5569_o = n5367_o[4]; // extract
  assign n5570_o = n5373_o[4]; // extract
  assign n5572_o = n5446_o[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5576_o = n5572_o;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5576_o = n5570_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5576_o = n5569_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5576_o = n5568_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5576_o = n5567_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5576_o = n5566_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5576_o = n5565_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5576_o = n5564_o;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5576_o = n5563_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5576_o = n5562_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5576_o = n5561_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5576_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5576_o = 1'b0;
      default: n5576_o = 1'b0;
    endcase
  assign n5577_o = n5229_o[5]; // extract
  assign n5578_o = n5236_o[5]; // extract
  assign n5579_o = n5241_o[5]; // extract
  assign n5580_o = n5248_o[5]; // extract
  assign n5581_o = n5257_o[5]; // extract
  assign n5582_o = n5290_o[5]; // extract
  assign n5583_o = n5296_o[5]; // extract
  assign n5584_o = n5367_o[5]; // extract
  assign n5585_o = n5373_o[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5590_o = n5585_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5590_o = n5584_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5590_o = n5583_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5590_o = n5582_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5590_o = n5581_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5590_o = n5580_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5590_o = n5579_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5590_o = n5578_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5590_o = n5577_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5590_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5590_o = 1'b0;
      default: n5590_o = 1'b0;
    endcase
  assign n5591_o = n5229_o[6]; // extract
  assign n5592_o = n5236_o[6]; // extract
  assign n5593_o = n5241_o[6]; // extract
  assign n5594_o = n5248_o[6]; // extract
  assign n5595_o = n5257_o[6]; // extract
  assign n5596_o = n5290_o[6]; // extract
  assign n5597_o = n5296_o[6]; // extract
  assign n5598_o = n5367_o[6]; // extract
  assign n5599_o = n5373_o[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5604_o = n5599_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5604_o = n5598_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5604_o = n5597_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5604_o = n5596_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5604_o = n5595_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5604_o = n5594_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5604_o = n5593_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5604_o = n5592_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5604_o = n5591_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5604_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5604_o = 1'b0;
      default: n5604_o = 1'b0;
    endcase
  assign n5605_o = n5229_o[7]; // extract
  assign n5606_o = n5236_o[7]; // extract
  assign n5607_o = n5241_o[7]; // extract
  assign n5608_o = n5248_o[7]; // extract
  assign n5609_o = n5257_o[7]; // extract
  assign n5610_o = n5290_o[7]; // extract
  assign n5611_o = n5296_o[7]; // extract
  assign n5612_o = n5367_o[7]; // extract
  assign n5613_o = n5373_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b1;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5618_o = n5613_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5618_o = n5612_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5618_o = n5611_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5618_o = n5610_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5618_o = n5609_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5618_o = n5252_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5618_o = n5608_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5618_o = n5607_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5618_o = n5606_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5618_o = n5605_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5618_o = n5224_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5618_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5618_o = n5194_o;
      default: n5618_o = 1'b0;
    endcase
  assign n5619_o = n5229_o[8]; // extract
  assign n5620_o = n5236_o[8]; // extract
  assign n5621_o = n5241_o[8]; // extract
  assign n5622_o = n5248_o[8]; // extract
  assign n5623_o = n5257_o[8]; // extract
  assign n5624_o = n5290_o[8]; // extract
  assign n5625_o = n5296_o[8]; // extract
  assign n5626_o = n5367_o[8]; // extract
  assign n5627_o = n5373_o[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5632_o = 1'b1;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5632_o = n5627_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5632_o = n5626_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5632_o = n5625_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5632_o = n5624_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5632_o = n5623_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5632_o = n5622_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5632_o = n5621_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5632_o = n5620_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5632_o = n5619_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5632_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5632_o = 1'b1;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5632_o = 1'b0;
      default: n5632_o = 1'b0;
    endcase
  assign n5633_o = n5229_o[9]; // extract
  assign n5634_o = n5236_o[9]; // extract
  assign n5635_o = n5241_o[9]; // extract
  assign n5636_o = n5248_o[9]; // extract
  assign n5637_o = n5257_o[9]; // extract
  assign n5638_o = n5290_o[9]; // extract
  assign n5639_o = n5296_o[9]; // extract
  assign n5640_o = n5367_o[9]; // extract
  assign n5641_o = n5373_o[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5646_o = 1'b1;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5646_o = n5641_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5646_o = n5640_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5646_o = n5639_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5646_o = n5638_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5646_o = n5637_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5646_o = n5636_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5646_o = n5635_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5646_o = n5634_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5646_o = n5633_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5646_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5646_o = 1'b0;
      default: n5646_o = 1'b0;
    endcase
  assign n5647_o = n5229_o[10]; // extract
  assign n5648_o = n5236_o[10]; // extract
  assign n5649_o = n5241_o[10]; // extract
  assign n5650_o = n5248_o[10]; // extract
  assign n5651_o = n5257_o[10]; // extract
  assign n5652_o = n5290_o[10]; // extract
  assign n5653_o = n5296_o[10]; // extract
  assign n5654_o = n5367_o[10]; // extract
  assign n5655_o = n5373_o[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5660_o = 1'b1;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5660_o = n5655_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5660_o = n5654_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5660_o = n5653_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5660_o = n5652_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5660_o = n5651_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5660_o = n5650_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5660_o = n5649_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5660_o = n5648_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5660_o = n5647_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5660_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5660_o = 1'b0;
      default: n5660_o = 1'b0;
    endcase
  assign n5661_o = n5197_o[0]; // extract
  assign n5662_o = n5229_o[11]; // extract
  assign n5663_o = n5236_o[11]; // extract
  assign n5664_o = n5241_o[11]; // extract
  assign n5665_o = n5248_o[11]; // extract
  assign n5666_o = n5257_o[11]; // extract
  assign n5667_o = n5290_o[11]; // extract
  assign n5668_o = n5296_o[11]; // extract
  assign n5669_o = n5367_o[11]; // extract
  assign n5670_o = n5373_o[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5675_o = n5670_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5675_o = n5669_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5675_o = n5668_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5675_o = n5667_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5675_o = n5666_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5675_o = n5253_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5675_o = n5665_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5675_o = n5664_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5675_o = n5663_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5675_o = n5662_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5675_o = n5225_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5675_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5675_o = n5661_o;
      default: n5675_o = 1'b0;
    endcase
  assign n5676_o = n5197_o[1]; // extract
  assign n5677_o = n5229_o[12]; // extract
  assign n5678_o = n5236_o[12]; // extract
  assign n5679_o = n5241_o[12]; // extract
  assign n5680_o = n5248_o[12]; // extract
  assign n5681_o = n5257_o[12]; // extract
  assign n5682_o = n5290_o[12]; // extract
  assign n5683_o = n5296_o[12]; // extract
  assign n5684_o = n5367_o[12]; // extract
  assign n5685_o = n5373_o[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5690_o = n5685_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5690_o = n5684_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5690_o = n5683_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5690_o = n5682_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5690_o = n5681_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5690_o = n5680_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5690_o = n5679_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5690_o = n5678_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5690_o = n5677_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5690_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5690_o = 1'b1;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5690_o = n5676_o;
      default: n5690_o = 1'b0;
    endcase
  assign n5691_o = n5229_o[15:13]; // extract
  assign n5692_o = n5236_o[15:13]; // extract
  assign n5693_o = n5241_o[15:13]; // extract
  assign n5694_o = n5248_o[15:13]; // extract
  assign n5695_o = n5257_o[15:13]; // extract
  assign n5696_o = n5290_o[15:13]; // extract
  assign n5697_o = n5296_o[15:13]; // extract
  assign n5698_o = n5367_o[15:13]; // extract
  assign n5699_o = n5373_o[15:13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5704_o = n5699_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5704_o = n5698_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5704_o = n5697_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5704_o = n5696_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5704_o = n5695_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5704_o = n5694_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5704_o = n5693_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5704_o = n5692_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5704_o = n5691_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5704_o = 3'b000;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5704_o = 3'b000;
      default: n5704_o = 3'b000;
    endcase
  assign n5705_o = n5226_o[0]; // extract
  assign n5706_o = n5229_o[16]; // extract
  assign n5707_o = n5236_o[16]; // extract
  assign n5708_o = n5241_o[16]; // extract
  assign n5709_o = n5248_o[16]; // extract
  assign n5710_o = n5254_o[0]; // extract
  assign n5711_o = n5257_o[16]; // extract
  assign n5712_o = n5290_o[16]; // extract
  assign n5713_o = n5296_o[16]; // extract
  assign n5714_o = n5367_o[16]; // extract
  assign n5715_o = n5373_o[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5720_o = 1'b1;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5720_o = n5715_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5720_o = n5714_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5720_o = n5713_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5720_o = n5712_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5720_o = n5711_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5720_o = n5710_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5720_o = n5709_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5720_o = n5708_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5720_o = n5707_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5720_o = n5706_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5720_o = n5705_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5720_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5720_o = 1'b0;
      default: n5720_o = 1'b0;
    endcase
  assign n5721_o = n5226_o[1]; // extract
  assign n5722_o = n5229_o[17]; // extract
  assign n5723_o = n5236_o[17]; // extract
  assign n5724_o = n5241_o[17]; // extract
  assign n5725_o = n5248_o[17]; // extract
  assign n5726_o = n5254_o[1]; // extract
  assign n5727_o = n5257_o[17]; // extract
  assign n5728_o = n5290_o[17]; // extract
  assign n5729_o = n5296_o[17]; // extract
  assign n5730_o = n5367_o[17]; // extract
  assign n5731_o = n5373_o[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5736_o = n5731_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5736_o = n5730_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5736_o = n5729_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5736_o = n5728_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5736_o = n5727_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5736_o = n5726_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5736_o = n5725_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5736_o = n5724_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5736_o = n5723_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5736_o = n5722_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5736_o = n5721_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5736_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5736_o = n5198_o;
      default: n5736_o = 1'b0;
    endcase
  assign n5737_o = n5226_o[3:2]; // extract
  assign n5738_o = n5229_o[19:18]; // extract
  assign n5739_o = n5236_o[19:18]; // extract
  assign n5740_o = n5241_o[19:18]; // extract
  assign n5741_o = n5248_o[19:18]; // extract
  assign n5742_o = n5254_o[3:2]; // extract
  assign n5743_o = n5257_o[19:18]; // extract
  assign n5744_o = n5290_o[19:18]; // extract
  assign n5745_o = n5296_o[19:18]; // extract
  assign n5746_o = n5367_o[19:18]; // extract
  assign n5747_o = n5373_o[19:18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5752_o = 2'b10;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5752_o = n5747_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5752_o = n5746_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5752_o = n5745_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5752_o = n5744_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5752_o = n5743_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5752_o = n5742_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5752_o = n5741_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5752_o = n5740_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5752_o = n5739_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5752_o = n5738_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5752_o = n5737_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5752_o = 2'b00;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5752_o = 2'b00;
      default: n5752_o = 2'b00;
    endcase
  assign n5753_o = n5226_o[4]; // extract
  assign n5754_o = n5229_o[20]; // extract
  assign n5755_o = n5236_o[20]; // extract
  assign n5756_o = n5241_o[20]; // extract
  assign n5757_o = n5248_o[20]; // extract
  assign n5758_o = n5254_o[4]; // extract
  assign n5759_o = n5257_o[20]; // extract
  assign n5760_o = n5290_o[20]; // extract
  assign n5761_o = n5296_o[20]; // extract
  assign n5762_o = n5367_o[20]; // extract
  assign n5763_o = n5373_o[20]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5768_o = n5763_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5768_o = n5762_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5768_o = n5761_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5768_o = n5760_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5768_o = n5759_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5768_o = n5758_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5768_o = n5757_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5768_o = n5756_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5768_o = n5755_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5768_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5768_o = n5754_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5768_o = n5753_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5768_o = 1'b1;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5768_o = 1'b0;
      default: n5768_o = 1'b0;
    endcase
  assign n5769_o = n5226_o[5]; // extract
  assign n5770_o = n5229_o[21]; // extract
  assign n5771_o = n5236_o[21]; // extract
  assign n5772_o = n5241_o[21]; // extract
  assign n5773_o = n5248_o[21]; // extract
  assign n5774_o = n5254_o[5]; // extract
  assign n5775_o = n5257_o[21]; // extract
  assign n5776_o = n5290_o[21]; // extract
  assign n5777_o = n5296_o[21]; // extract
  assign n5778_o = n5367_o[21]; // extract
  assign n5779_o = n5373_o[21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5784_o = n5779_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5784_o = n5778_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5784_o = n5777_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5784_o = n5776_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5784_o = n5775_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5784_o = n5774_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5784_o = n5773_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5784_o = n5772_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5784_o = n5771_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5784_o = n5770_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5784_o = n5769_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5784_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5784_o = n5202_o;
      default: n5784_o = 1'b0;
    endcase
  assign n5785_o = n5226_o[6]; // extract
  assign n5786_o = n5229_o[22]; // extract
  assign n5787_o = n5236_o[22]; // extract
  assign n5788_o = n5241_o[22]; // extract
  assign n5789_o = n5248_o[22]; // extract
  assign n5790_o = n5254_o[6]; // extract
  assign n5791_o = n5257_o[22]; // extract
  assign n5792_o = n5290_o[22]; // extract
  assign n5793_o = n5296_o[22]; // extract
  assign n5794_o = n5367_o[22]; // extract
  assign n5795_o = n5373_o[22]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5800_o = n5795_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5800_o = n5794_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5800_o = n5793_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5800_o = n5792_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5800_o = n5791_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5800_o = n5790_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5800_o = n5789_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5800_o = n5788_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5800_o = n5787_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5800_o = n5786_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5800_o = n5785_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5800_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5800_o = 1'b0;
      default: n5800_o = 1'b0;
    endcase
  assign n5801_o = n5226_o[7]; // extract
  assign n5802_o = n5229_o[23]; // extract
  assign n5803_o = n5236_o[23]; // extract
  assign n5804_o = n5241_o[23]; // extract
  assign n5805_o = n5248_o[23]; // extract
  assign n5806_o = n5254_o[7]; // extract
  assign n5807_o = n5257_o[23]; // extract
  assign n5808_o = n5290_o[23]; // extract
  assign n5809_o = n5296_o[23]; // extract
  assign n5810_o = n5367_o[23]; // extract
  assign n5811_o = n5373_o[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5816_o = n5811_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5816_o = n5810_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5816_o = n5809_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5816_o = n5808_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5816_o = n5807_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5816_o = n5806_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5816_o = n5805_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5816_o = n5804_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5816_o = n5803_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5816_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5816_o = n5802_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5816_o = n5801_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5816_o = 1'b1;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5816_o = 1'b0;
      default: n5816_o = 1'b0;
    endcase
  assign n5817_o = n5226_o[12:8]; // extract
  assign n5818_o = n5229_o[28:24]; // extract
  assign n5819_o = n5236_o[28:24]; // extract
  assign n5820_o = n5241_o[28:24]; // extract
  assign n5821_o = n5248_o[28:24]; // extract
  assign n5822_o = n5254_o[12:8]; // extract
  assign n5823_o = n5257_o[28:24]; // extract
  assign n5824_o = n5290_o[28:24]; // extract
  assign n5825_o = n5296_o[28:24]; // extract
  assign n5826_o = n5367_o[28:24]; // extract
  assign n5827_o = n5373_o[28:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00001;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5832_o = n5827_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5832_o = n5826_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5832_o = n5825_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5832_o = n5824_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5832_o = n5823_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5832_o = n5822_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5832_o = n5821_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5832_o = n5820_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5832_o = n5819_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5832_o = n5818_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5832_o = n5817_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5832_o = 5'b00000;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5832_o = 5'b00000;
      default: n5832_o = 5'b00000;
    endcase
  assign n5833_o = n5226_o[13]; // extract
  assign n5834_o = n5229_o[29]; // extract
  assign n5835_o = n5236_o[29]; // extract
  assign n5836_o = n5241_o[29]; // extract
  assign n5837_o = n5248_o[29]; // extract
  assign n5838_o = n5254_o[13]; // extract
  assign n5839_o = n5257_o[29]; // extract
  assign n5840_o = n5290_o[29]; // extract
  assign n5841_o = n5296_o[29]; // extract
  assign n5842_o = n5367_o[29]; // extract
  assign n5843_o = n5373_o[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5848_o = n5843_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5848_o = n5842_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5848_o = n5841_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5848_o = n5840_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5848_o = n5839_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5848_o = n5838_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5848_o = n5837_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5848_o = n5836_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5848_o = n5835_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5848_o = n5834_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5848_o = n5833_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5848_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5848_o = 1'b0;
      default: n5848_o = 1'b0;
    endcase
  assign n5849_o = n5220_o[0]; // extract
  assign n5850_o = n5226_o[14]; // extract
  assign n5851_o = n5229_o[30]; // extract
  assign n5852_o = n5236_o[30]; // extract
  assign n5853_o = n5241_o[30]; // extract
  assign n5854_o = n5248_o[30]; // extract
  assign n5855_o = n5254_o[14]; // extract
  assign n5856_o = n5257_o[30]; // extract
  assign n5857_o = n5290_o[30]; // extract
  assign n5858_o = n5296_o[30]; // extract
  assign n5859_o = n5367_o[30]; // extract
  assign n5860_o = n5373_o[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b1;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5865_o = n5860_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5865_o = n5859_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5865_o = n5858_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5865_o = n5857_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5865_o = n5856_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5865_o = n5855_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5865_o = n5854_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5865_o = n5853_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5865_o = n5852_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5865_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5865_o = n5851_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5865_o = n5850_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5865_o = n5849_o;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5865_o = 1'b0;
      default: n5865_o = 1'b0;
    endcase
  assign n5866_o = n5220_o[1]; // extract
  assign n5867_o = n5226_o[15]; // extract
  assign n5868_o = n5229_o[31]; // extract
  assign n5869_o = n5236_o[31]; // extract
  assign n5870_o = n5241_o[31]; // extract
  assign n5871_o = n5248_o[31]; // extract
  assign n5872_o = n5254_o[15]; // extract
  assign n5873_o = n5257_o[31]; // extract
  assign n5874_o = n5290_o[31]; // extract
  assign n5875_o = n5296_o[31]; // extract
  assign n5876_o = n5367_o[31]; // extract
  assign n5877_o = n5373_o[31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1936:5  */
  always @*
    case (n5496_o)
      66'b100000000000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b1;
      66'b010000000000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b001000000000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000100000000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000010000000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000001000000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000100000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000010000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000001000000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000100000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000010000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000001000000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000100000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000010000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000001000000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000100000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000010000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000001000000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000100000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000010000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000001000000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000100000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000010000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000001000000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000100000000000000000000000000000000000000000: n5882_o = n5877_o;
      66'b000000000000000000000000010000000000000000000000000000000000000000: n5882_o = n5876_o;
      66'b000000000000000000000000001000000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000100000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000010000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000001000000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000100000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000010000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000001000000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000100000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000010000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000001000000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000100000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000010000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000001000000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000100000000000000000000000000: n5882_o = n5875_o;
      66'b000000000000000000000000000000000000000010000000000000000000000000: n5882_o = n5874_o;
      66'b000000000000000000000000000000000000000001000000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000100000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000010000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000001000000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000100000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000010000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000001000000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000100000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000010000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000001000000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000100000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000010000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000001000000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000100000000000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000010000000000: n5882_o = n5873_o;
      66'b000000000000000000000000000000000000000000000000000000001000000000: n5882_o = n5872_o;
      66'b000000000000000000000000000000000000000000000000000000000100000000: n5882_o = n5871_o;
      66'b000000000000000000000000000000000000000000000000000000000010000000: n5882_o = n5244_o;
      66'b000000000000000000000000000000000000000000000000000000000001000000: n5882_o = n5870_o;
      66'b000000000000000000000000000000000000000000000000000000000000100000: n5882_o = n5869_o;
      66'b000000000000000000000000000000000000000000000000000000000000010000: n5882_o = 1'b0;
      66'b000000000000000000000000000000000000000000000000000000000000001000: n5882_o = n5868_o;
      66'b000000000000000000000000000000000000000000000000000000000000000100: n5882_o = n5867_o;
      66'b000000000000000000000000000000000000000000000000000000000000000010: n5882_o = n5866_o;
      66'b000000000000000000000000000000000000000000000000000000000000000001: n5882_o = 1'b0;
      default: n5882_o = 1'b0;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2143:16  */
  assign n5910_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2147:21  */
  assign n5914_o = csr[30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2148:15  */
  assign n5915_o = csr[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2149:32  */
  assign n5916_o = csr_rdata | xcsr_rdata;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2148:7  */
  assign n5918_o = n5915_o ? n5916_o : 32'b00000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2157:22  */
  assign n5926_o = csr[94:63]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2172:13  */
  assign n5930_o = csr[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2172:36  */
  assign n5931_o = csr[11:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2172:50  */
  assign n5933_o = n5931_o == 4'b1011;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2172:23  */
  assign n5934_o = n5933_o & n5930_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2173:19  */
  assign n5935_o = csr[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2173:23  */
  assign n5936_o = ~n5935_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:47  */
  assign n5937_o = csr[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:47  */
  assign n5942_o = csr[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2173:7  */
  assign n5947_o = n5936_o ? n6362_o : 16'b0000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2173:7  */
  assign n5948_o = n5936_o ? 16'b0000000000000000 : n6431_o;
  assign n5949_o = {n5948_o, n5947_o};
  assign n5950_o = {16'b0000000000000000, 16'b0000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2172:5  */
  assign n5951_o = n5934_o ? n5949_o : n5950_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:18  */
  assign n5954_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2195:22  */
  assign n5959_o = cnt[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2196:28  */
  assign n5960_o = csr[62:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2198:34  */
  assign n5961_o = cnt[337:306]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2195:9  */
  assign n5962_o = n5959_o ? n5960_o : n5961_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2200:36  */
  assign n5963_o = cnt[338]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2202:22  */
  assign n5964_o = cnt[16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2203:28  */
  assign n5965_o = csr[62:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:57  */
  assign n5966_o = cnt[239:208]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:80  */
  assign n5967_o = cnt[341]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:62  */
  assign n5968_o = {31'b0, n5967_o};  //  uext
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:62  */
  assign n5969_o = n5966_o + n5968_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2202:9  */
  assign n5970_o = n5964_o ? n5965_o : n5969_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:58  */
  assign n5981_o = cnt[143:112]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:50  */
  assign n5983_o = {1'b0, n5981_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:63  */
  assign n5985_o = n5983_o + 33'b000000000000000000000000000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:81  */
  assign n5986_o = cnt[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:68  */
  assign n5987_o = n5986_o ? n5985_o : n5992_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:58  */
  assign n5988_o = cnt[143:112]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:50  */
  assign n5990_o = {1'b0, n5988_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:63  */
  assign n5992_o = n5990_o + 33'b000000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:18  */
  assign n5994_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2195:22  */
  assign n5999_o = cnt[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2196:28  */
  assign n6000_o = csr[62:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2198:34  */
  assign n6001_o = cnt[304:273]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2195:9  */
  assign n6002_o = n5999_o ? n6000_o : n6001_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2200:36  */
  assign n6003_o = cnt[305]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2202:22  */
  assign n6004_o = cnt[17]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2203:28  */
  assign n6005_o = csr[62:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:57  */
  assign n6006_o = cnt[207:176]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:80  */
  assign n6007_o = cnt[340]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:62  */
  assign n6008_o = {31'b0, n6007_o};  //  uext
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:62  */
  assign n6009_o = n6006_o + n6008_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2202:9  */
  assign n6010_o = n6004_o ? n6005_o : n6009_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:58  */
  assign n6021_o = cnt[111:80]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:50  */
  assign n6023_o = {1'b0, n6021_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:63  */
  assign n6025_o = n6023_o + 33'b000000000000000000000000000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:81  */
  assign n6026_o = cnt[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:68  */
  assign n6027_o = n6026_o ? n6025_o : n6032_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:58  */
  assign n6028_o = cnt[111:80]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:50  */
  assign n6030_o = {1'b0, n6028_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:63  */
  assign n6032_o = n6030_o + 33'b000000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:18  */
  assign n6034_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2195:22  */
  assign n6039_o = cnt[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2196:28  */
  assign n6040_o = csr[62:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2198:34  */
  assign n6041_o = cnt[271:240]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2195:9  */
  assign n6042_o = n6039_o ? n6040_o : n6041_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2200:36  */
  assign n6043_o = cnt[272]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2202:22  */
  assign n6044_o = cnt[18]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2203:28  */
  assign n6045_o = csr[62:31]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:57  */
  assign n6046_o = cnt[175:144]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:80  */
  assign n6047_o = cnt[339]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:62  */
  assign n6048_o = {31'b0, n6047_o};  //  uext
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2205:62  */
  assign n6049_o = n6046_o + n6048_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2202:9  */
  assign n6050_o = n6044_o ? n6045_o : n6049_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:58  */
  assign n6061_o = cnt[79:48]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:50  */
  assign n6063_o = {1'b0, n6061_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:63  */
  assign n6065_o = n6063_o + 33'b000000000000000000000000000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:81  */
  assign n6066_o = cnt[34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2211:68  */
  assign n6067_o = n6066_o ? n6065_o : n6072_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:58  */
  assign n6068_o = cnt[79:48]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:50  */
  assign n6070_o = {1'b0, n6068_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2212:63  */
  assign n6072_o = n6070_o + 33'b000000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2224:29  */
  assign n6074_o = cnt[143:112]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2225:29  */
  assign n6077_o = cnt[239:208]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2226:29  */
  assign n6080_o = cnt[79:48]; // extract
  assign n6081_o = n6075_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2227:29  */
  assign n6082_o = cnt[175:144]; // extract
  assign n6083_o = n6078_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2299:16  */
  assign n6088_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2305:32  */
  assign n6092_o = cnt_event[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2305:78  */
  assign n6093_o = csr[321]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2305:57  */
  assign n6094_o = ~n6093_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2305:52  */
  assign n6095_o = n6092_o & n6094_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2305:103  */
  assign n6096_o = debug_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2305:88  */
  assign n6097_o = ~n6096_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2305:83  */
  assign n6098_o = n6095_o & n6097_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2306:32  */
  assign n6100_o = cnt_event[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2306:78  */
  assign n6101_o = csr[323]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2306:57  */
  assign n6102_o = ~n6101_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2306:52  */
  assign n6103_o = n6100_o & n6102_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2306:103  */
  assign n6104_o = debug_ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2306:88  */
  assign n6105_o = ~n6104_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2306:83  */
  assign n6106_o = n6103_o & n6105_o;
  assign n6107_o = n6091_o[15:3]; // extract
  assign n6108_o = n6091_o[1]; // extract
  assign n6109_o = {n6107_o, n6106_o, n6108_o, n6098_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2318:56  */
  assign n6115_o = ~sleep_mode;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2318:39  */
  assign n6116_o = n6115_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2320:60  */
  assign n6120_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2320:66  */
  assign n6122_o = n6120_o == 4'b0110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2320:39  */
  assign n6123_o = n6122_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2323:66  */
  assign n6126_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2323:72  */
  assign n6128_o = n6126_o == 4'b0110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2323:104  */
  assign n6129_o = execute_engine[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2323:84  */
  assign n6130_o = n6129_o & n6128_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2323:45  */
  assign n6131_o = n6130_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2324:66  */
  assign n6134_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2324:72  */
  assign n6136_o = n6134_o == 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2324:102  */
  assign n6137_o = issue_engine[86:85]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2324:110  */
  assign n6139_o = n6137_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2324:84  */
  assign n6140_o = n6139_o & n6136_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2324:45  */
  assign n6141_o = n6140_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2325:66  */
  assign n6144_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2325:72  */
  assign n6146_o = n6144_o == 4'b0111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2325:45  */
  assign n6147_o = n6146_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2327:66  */
  assign n6150_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2327:72  */
  assign n6152_o = n6150_o == 4'b1000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2327:45  */
  assign n6153_o = n6152_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2328:66  */
  assign n6156_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2328:72  */
  assign n6158_o = n6156_o == 4'b1001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2328:45  */
  assign n6159_o = n6158_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2330:56  */
  assign n6162_o = ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2330:81  */
  assign n6163_o = ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2330:88  */
  assign n6164_o = ~n6163_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2330:71  */
  assign n6165_o = n6164_o & n6162_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2330:45  */
  assign n6166_o = n6165_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2331:56  */
  assign n6169_o = ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2331:81  */
  assign n6170_o = ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2331:71  */
  assign n6171_o = n6170_o & n6169_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2331:45  */
  assign n6172_o = n6171_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2332:56  */
  assign n6175_o = ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2332:64  */
  assign n6176_o = ~n6175_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2332:91  */
  assign n6177_o = execute_engine[3:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2332:97  */
  assign n6179_o = n6177_o == 4'b1100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2332:71  */
  assign n6180_o = n6179_o & n6176_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2332:45  */
  assign n6181_o = n6180_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2334:61  */
  assign n6184_o = trap_ctrl[95]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2334:45  */
  assign n6185_o = n6184_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2388:36  */
  assign n6194_o = csr[337]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2391:36  */
  assign n6197_o = csr[338]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2391:49  */
  assign n6199_o = 1'b1 ? n6197_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2395:36  */
  assign n6204_o = csr[343:341]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2399:36  */
  assign n6208_o = csr[339]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2400:47  */
  assign n6209_o = csr[340]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2400:47  */
  assign n6210_o = csr[340]; // extract
  assign n6211_o = {n6209_o, n6210_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2442:38  */
  assign n6215_o = csr[443]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2451:46  */
  assign n6223_o = csr[442]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2451:40  */
  assign n6225_o = {3'b000, n6223_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2458:38  */
  assign n6233_o = csr[441]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:358:5  */
  always @(posedge clk_i or posedge n2372_o)
    if (n2372_o)
      n6236_q <= 1'b1;
    else
      n6236_q <= n2430_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:358:5  */
  always @(posedge clk_i or posedge n2372_o)
    if (n2372_o)
      n6237_q <= n2436_o;
    else
      n6237_q <= n2431_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:353:5  */
  assign n6238_o = {n6236_q, n2458_o, n3326_o, n6237_q};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:353:5  */
  assign n6239_o = {prefetch_buffer_n2_prefetch_buffer_inst_avail_o, prefetch_buffer_n1_prefetch_buffer_inst_avail_o, prefetch_buffer_n2_prefetch_buffer_inst_free_o, prefetch_buffer_n1_prefetch_buffer_inst_free_o, n2618_o, n2615_o, n2486_o, n2478_o, prefetch_buffer_n1_prefetch_buffer_inst_rdata_o, prefetch_buffer_n2_prefetch_buffer_inst_rdata_o, n2462_o, n2466_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:491:7  */
  always @(posedge clk_i or posedge n2517_o)
    if (n2517_o)
      n6240_q <= 1'b0;
    else
      n6240_q <= n2531_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:489:7  */
  assign n6241_o = {n3327_o, n2611_o, neorv32_cpu_decompressor_inst_true_neorv32_cpu_decompressor_inst_ci_instr32_o, n2514_o, n2610_o, n2568_o, n6240_q};
  assign n6242_o = {n2958_o, n2952_o, 1'b0, 1'b0, 1'b0, n2946_o, 1'b0, 1'b0, 1'b0, n2962_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  assign n6243_o = execute_engine[203:172]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  assign n6244_o = n2821_o ? n2824_o : n6243_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  always @(posedge clk_i or posedge n2802_o)
    if (n2802_o)
      n6245_q <= 32'b00000000000000000000000000000000;
    else
      n6245_q <= n6244_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  always @(posedge clk_i or posedge n2802_o)
    if (n2802_o)
      n6246_q <= 32'b00000000000000000000000000000000;
    else
      n6246_q <= n2870_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  assign n6247_o = execute_engine[106:75]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  assign n6248_o = n2813_o ? n2816_o : n6247_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  always @(posedge clk_i or posedge n2802_o)
    if (n2802_o)
      n6249_q <= 32'b00000000000000000000000000000000;
    else
      n6249_q <= n6248_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  always @(posedge clk_i or posedge n2802_o)
    if (n2802_o)
      n6250_q <= 1'b0;
    else
      n6250_q <= n2812_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  always @(posedge clk_i or posedge n2802_o)
    if (n2802_o)
      n6251_q <= 32'b00000000000000000000000000000000;
    else
      n6251_q <= n2811_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  always @(posedge clk_i or posedge n2802_o)
    if (n2802_o)
      n6252_q <= 4'b0011;
    else
      n6252_q <= n2810_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:611:5  */
  assign n6253_o = {n6245_q, 28'b0000000000000000000000000000, n2913_o, n6246_q, n3331_o, n6249_q, n2799_o, n3330_o, n6250_q, n3329_o, n6251_q, n3328_o, n6252_q};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1138:5  */
  always @(posedge clk_i or posedge n3445_o)
    if (n3445_o)
      n6254_q <= 10'b0000000000;
    else
      n6254_q <= n3450_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1136:5  */
  assign n6255_o = {n3461_o, n3459_o, n6254_q};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1075:5  */
  always @(posedge clk_aux_i or posedge n3373_o)
    if (n3373_o)
      n6256_q <= 1'b0;
    else
      n6256_q <= n3387_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1551:5  */
  always @(posedge clk_i or posedge n4687_o)
    if (n4687_o)
      n6257_q <= 1'b0;
    else
      n6257_q <= n4706_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1502:5  */
  always @(posedge clk_i or posedge n4580_o)
    if (n4580_o)
      n6258_q <= 7'b0000000;
    else
      n6258_q <= n4681_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1442:5  */
  always @(posedge clk_aux_i or posedge n4272_o)
    if (n4272_o)
      n6259_q <= n4576_o;
    else
      n6259_q <= n4573_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1390:5  */
  always @(posedge clk_i or posedge n4206_o)
    if (n4206_o)
      n6260_q <= 11'b00000000000;
    else
      n6260_q <= n4266_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1388:5  */
  assign n6261_o = {1'b0, n3336_o, n4203_o, n2905_o, n3334_o, n4765_o, n3333_o, n3332_o, n6257_q, n4867_o, n6258_q, n4863_o, n6259_q, n4798_o, n6260_q};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:619:5  */
  always @(posedge clk_i or posedge n2802_o)
    if (n2802_o)
      n6262_q <= 67'b0000000000000000000000000000000000000000000000000000000000000000000;
    else
      n6262_q <= ctrl_nxt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:611:5  */
  assign n6263_o = {n3367_o, n3356_o, n3368_o, n3029_o, n3354_o, n3366_o, n3352_o, n3350_o, n3364_o, n3348_o, n3346_o, n2981_o, n3028_o, n2996_o, n3344_o, n3342_o, n3340_o, n3359_o, n3338_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2146:5  */
  always @(posedge clk_i or posedge n5910_o)
    if (n5910_o)
      n6264_q <= 32'b00000000000000000000000000000000;
    else
      n6264_q <= n5918_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2146:5  */
  always @(posedge clk_i or posedge n5910_o)
    if (n5910_o)
      n6265_q <= 1'b0;
    else
      n6265_q <= n5914_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1667:5  */
  always @(posedge clk_i or posedge n4910_o)
    if (n4910_o)
      n6266_q <= 32'b00000000000000000000000000000000;
    else
      n6266_q <= 32'b00000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1667:5  */
  always @(posedge clk_i or posedge n4910_o)
    if (n4910_o)
      n6267_q <= n5158_o;
    else
      n6267_q <= n5140_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1667:5  */
  always @(posedge clk_i or posedge n4910_o)
    if (n4910_o)
      n6268_q <= n5157_o;
    else
      n6268_q <= n5139_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1667:5  */
  always @(posedge clk_i or posedge n4910_o)
    if (n4910_o)
      n6269_q <= n5156_o;
    else
      n6269_q <= n5138_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1667:5  */
  always @(posedge clk_i or posedge n4910_o)
    if (n4910_o)
      n6270_q <= 1'b1;
    else
      n6270_q <= n5112_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1667:5  */
  always @(posedge clk_i or posedge n4910_o)
    if (n4910_o)
      n6271_q <= n5155_o;
    else
      n6271_q <= n5137_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1667:5  */
  always @(posedge clk_i or posedge n4910_o)
    if (n4910_o)
      n6272_q <= 1'b0;
    else
      n6272_q <= n4945_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1636:5  */
  assign n6273_o = {n6266_q, 4'b0110, n6215_o, 1'b0, 1'b0, 1'b0, 1'b0, hw_trigger_fired, 1'b0, 2'b00, 3'b000, n6225_o, 1'b0, 4'b0000, 1'b1, 1'b0, 1'b0, 1'b1, n6233_o, 1'b0, 1'b0, n6267_q, n5185_o, n6268_q, 4'b0100, 12'b000000000000, n6194_o, 1'b0, 1'b0, n6199_o, 1'b0, 1'b1, 1'b0, n6204_o, 1'b0, 1'b1, 1'b0, n6208_o, n6211_o, n6269_q, n5189_o, n6270_q, n5175_o, n6271_q, n4890_o, n6264_q, n4905_o, n3370_o, n6265_q, n3369_o, n6272_q, n4877_o, n4876_o, n4869_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2301:5  */
  always @(posedge clk_i or posedge n6088_o)
    if (n6088_o)
      n6275_q <= 16'b0000000000000000;
    else
      n6275_q <= n6109_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n6034_o)
    if (n6034_o)
      n6276_q <= 1'b0;
    else
      n6276_q <= n6043_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n6034_o)
    if (n6034_o)
      n6277_q <= 32'b00000000000000000000000000000000;
    else
      n6277_q <= n6050_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n6034_o)
    if (n6034_o)
      n6278_q <= 32'b00000000000000000000000000000000;
    else
      n6278_q <= n6042_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n5994_o)
    if (n5994_o)
      n6279_q <= 1'b0;
    else
      n6279_q <= n6003_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n5994_o)
    if (n5994_o)
      n6280_q <= 32'b00000000000000000000000000000000;
    else
      n6280_q <= n6010_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n5994_o)
    if (n5994_o)
      n6281_q <= 32'b00000000000000000000000000000000;
    else
      n6281_q <= n6002_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n5954_o)
    if (n5954_o)
      n6282_q <= 1'b0;
    else
      n6282_q <= n5963_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n5954_o)
    if (n5954_o)
      n6283_q <= 32'b00000000000000000000000000000000;
    else
      n6283_q <= n5970_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2193:7  */
  always @(posedge clk_i or posedge n5954_o)
    if (n5954_o)
      n6284_q <= 32'b00000000000000000000000000000000;
    else
      n6284_q <= n5962_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:7  */
  assign n6285_o = {n6282_q, n6279_q, n6276_q, n5987_o, n6027_o, n6067_o, n6283_q, n6280_q, n6277_q, n6284_q, n6281_q, n6278_q, n6275_q, n5951_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:7  */
  assign n6286_o = {n6074_o, n6081_o, n6080_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:7  */
  assign n6287_o = {n6077_o, n6083_o, n6082_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:7  */
  assign n6288_o = {n6185_o, n6181_o, n6172_o, n6166_o, n6159_o, n6153_o, n6147_o, n6141_o, n6131_o, n6123_o, 1'b0, n6116_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:7  */
  assign n6289_o = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:7  */
  assign n6290_o = {n5882_o, n5865_o, n5848_o, n5832_o, n5816_o, n5800_o, n5784_o, n5768_o, n5752_o, n5736_o, n5720_o, n5704_o, n5690_o, n5675_o, n5660_o, n5646_o, n5632_o, n5618_o, n5604_o, n5590_o, n5576_o, n5560_o, n5544_o, n5528_o, n5512_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:7  */
  assign n6291_o = {n3443_o, n3442_o, sleep_mode, n3441_o, n3440_o, n3439_o, n3438_o, n3436_o, n3433_o, n3431_o, n3426_o, n3425_o, n3424_o, n3423_o, n3422_o, n3421_o, n3420_o, n3419_o, n3418_o, n3417_o, n3416_o, n3415_o, n3414_o, n3413_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2189:7  */
  assign n6292_o = {n2494_o, 1'b0, n2488_o, 1'b1, 1'b0, n2454_o, 4'b0000, 32'b00000000000000000000000000000000, n2442_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:552:5  */
  always @(posedge clk_i or posedge n2620_o)
    if (n2620_o)
      n6293_q <= 32'b00000000000000000000000000000000;
    else
      n6293_q <= n2781_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6294_o = n5937_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6295_o = ~n6294_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6296_o = n5937_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6297_o = ~n6296_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6298_o = n6295_o & n6297_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6299_o = n6295_o & n6296_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6300_o = n6294_o & n6297_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6301_o = n6294_o & n6296_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6302_o = n5937_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6303_o = ~n6302_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6304_o = n6298_o & n6303_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6305_o = n6298_o & n6302_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6306_o = n6299_o & n6303_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6307_o = n6299_o & n6302_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6308_o = n6300_o & n6303_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6309_o = n6300_o & n6302_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6310_o = n6301_o & n6303_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6311_o = n6301_o & n6302_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6312_o = n5937_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6313_o = ~n6312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6314_o = n6304_o & n6313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6315_o = n6304_o & n6312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6316_o = n6305_o & n6313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6317_o = n6305_o & n6312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6318_o = n6306_o & n6313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6319_o = n6306_o & n6312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6320_o = n6307_o & n6313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6321_o = n6307_o & n6312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6322_o = n6308_o & n6313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6323_o = n6308_o & n6312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6324_o = n6309_o & n6313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6325_o = n6309_o & n6312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6326_o = n6310_o & n6313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6327_o = n6310_o & n6312_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6328_o = n6311_o & n6313_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6329_o = n6311_o & n6312_o;
  assign n6330_o = n5928_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6331_o = n6314_o ? 1'b1 : n6330_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2187:5  */
  assign n6332_o = n5928_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6333_o = n6315_o ? 1'b1 : n6332_o;
  assign n6334_o = n5928_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6335_o = n6316_o ? 1'b1 : n6334_o;
  assign n6336_o = n5928_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6337_o = n6317_o ? 1'b1 : n6336_o;
  assign n6338_o = n5928_o[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6339_o = n6318_o ? 1'b1 : n6338_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:19  */
  assign n6340_o = n5928_o[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6341_o = n6319_o ? 1'b1 : n6340_o;
  assign n6342_o = n5928_o[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6343_o = n6320_o ? 1'b1 : n6342_o;
  assign n6344_o = n5928_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6345_o = n6321_o ? 1'b1 : n6344_o;
  assign n6346_o = n5928_o[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6347_o = n6322_o ? 1'b1 : n6346_o;
  assign n6348_o = n5928_o[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6349_o = n6323_o ? 1'b1 : n6348_o;
  assign n6350_o = n5928_o[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6351_o = n6324_o ? 1'b1 : n6350_o;
  assign n6352_o = n5928_o[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6353_o = n6325_o ? 1'b1 : n6352_o;
  assign n6354_o = n5928_o[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6355_o = n6326_o ? 1'b1 : n6354_o;
  assign n6356_o = n5928_o[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6357_o = n6327_o ? 1'b1 : n6356_o;
  assign n6358_o = n5928_o[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6359_o = n6328_o ? 1'b1 : n6358_o;
  assign n6360_o = n5928_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2174:9  */
  assign n6361_o = n6329_o ? 1'b1 : n6360_o;
  assign n6362_o = {n6361_o, n6359_o, n6357_o, n6355_o, n6353_o, n6351_o, n6349_o, n6347_o, n6345_o, n6343_o, n6341_o, n6339_o, n6337_o, n6335_o, n6333_o, n6331_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6363_o = n5942_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6364_o = ~n6363_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6365_o = n5942_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6366_o = ~n6365_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6367_o = n6364_o & n6366_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6368_o = n6364_o & n6365_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6369_o = n6363_o & n6366_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6370_o = n6363_o & n6365_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6371_o = n5942_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6372_o = ~n6371_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6373_o = n6367_o & n6372_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6374_o = n6367_o & n6371_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6375_o = n6368_o & n6372_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6376_o = n6368_o & n6371_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6377_o = n6369_o & n6372_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6378_o = n6369_o & n6371_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6379_o = n6370_o & n6372_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6380_o = n6370_o & n6371_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6381_o = n5942_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6382_o = ~n6381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6383_o = n6373_o & n6382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6384_o = n6373_o & n6381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6385_o = n6374_o & n6382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6386_o = n6374_o & n6381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6387_o = n6375_o & n6382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6388_o = n6375_o & n6381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6389_o = n6376_o & n6382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6390_o = n6376_o & n6381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6391_o = n6377_o & n6382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6392_o = n6377_o & n6381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6393_o = n6378_o & n6382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6394_o = n6378_o & n6381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6395_o = n6379_o & n6382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6396_o = n6379_o & n6381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6397_o = n6380_o & n6382_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6398_o = n6380_o & n6381_o;
  assign n6399_o = n5929_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6400_o = n6383_o ? 1'b1 : n6399_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:716:12  */
  assign n6401_o = n5929_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6402_o = n6384_o ? 1'b1 : n6401_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:716:12  */
  assign n6403_o = n5929_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6404_o = n6385_o ? 1'b1 : n6403_o;
  assign n6405_o = n5929_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6406_o = n6386_o ? 1'b1 : n6405_o;
  assign n6407_o = n5929_o[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6408_o = n6387_o ? 1'b1 : n6407_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:716:12  */
  assign n6409_o = n5929_o[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6410_o = n6388_o ? 1'b1 : n6409_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:716:12  */
  assign n6411_o = n5929_o[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6412_o = n6389_o ? 1'b1 : n6411_o;
  assign n6413_o = n5929_o[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6414_o = n6390_o ? 1'b1 : n6413_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1547:3  */
  assign n6415_o = n5929_o[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6416_o = n6391_o ? 1'b1 : n6415_o;
  assign n6417_o = n5929_o[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6418_o = n6392_o ? 1'b1 : n6417_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1498:3  */
  assign n6419_o = n5929_o[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6420_o = n6393_o ? 1'b1 : n6419_o;
  assign n6421_o = n5929_o[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6422_o = n6394_o ? 1'b1 : n6421_o;
  assign n6423_o = n5929_o[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6424_o = n6395_o ? 1'b1 : n6423_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1386:3  */
  assign n6425_o = n5929_o[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6426_o = n6396_o ? 1'b1 : n6425_o;
  assign n6427_o = n5929_o[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6428_o = n6397_o ? 1'b1 : n6427_o;
  assign n6429_o = n5929_o[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:2176:9  */
  assign n6430_o = n6398_o ? 1'b1 : n6429_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu_control.vhd:1241:72  */
  assign n6431_o = {n6430_o, n6428_o, n6426_o, n6424_o, n6422_o, n6420_o, n6418_o, n6416_o, n6414_o, n6412_o, n6410_o, n6408_o, n6406_o, n6404_o, n6402_o, n6400_o};
endmodule

module neorv32_sysinfo_0_16384_8192_4_4_64_4_64_32_32_8_256_ad514a383a71baac85f4c0ffc48c0bd10a15d22b
  (input  clk_i,
   input  rstn_i,
   input  [31:0] bus_req_i_addr,
   input  [31:0] bus_req_i_data,
   input  [3:0] bus_req_i_ben,
   input  bus_req_i_stb,
   input  bus_req_i_rw,
   input  bus_req_i_src,
   input  bus_req_i_priv,
   input  bus_req_i_rvso,
   input  bus_req_i_fence,
   output [31:0] bus_rsp_o_data,
   output bus_rsp_o_ack,
   output bus_rsp_o_err);
  wire [73:0] n2123_o;
  wire [31:0] n2125_o;
  wire n2126_o;
  wire n2127_o;
  wire [127:0] sysinfo;
  wire n2138_o;
  wire n2142_o;
  wire n2146_o;
  wire n2150_o;
  wire n2154_o;
  wire n2158_o;
  wire n2162_o;
  wire n2166_o;
  wire n2170_o;
  wire n2174_o;
  wire n2178_o;
  wire n2185_o;
  wire n2189_o;
  wire n2193_o;
  wire n2197_o;
  wire n2201_o;
  wire n2205_o;
  wire n2209_o;
  wire n2213_o;
  wire n2217_o;
  wire n2221_o;
  wire n2225_o;
  wire n2229_o;
  wire n2233_o;
  wire n2237_o;
  wire n2241_o;
  wire n2245_o;
  wire n2249_o;
  wire n2253_o;
  wire [3:0] n2258_o;
  wire [3:0] n2263_o;
  wire [3:0] n2268_o;
  wire [3:0] n2273_o;
  wire [3:0] n2277_o;
  wire [3:0] n2281_o;
  wire [3:0] n2285_o;
  wire [3:0] n2289_o;
  wire n2292_o;
  wire n2300_o;
  wire n2301_o;
  wire n2302_o;
  wire n2303_o;
  wire [1:0] n2305_o;
  wire [1:0] n2308_o;
  wire [32:0] n2311_o;
  wire [32:0] n2312_o;
  wire [32:0] n2313_o;
  wire [33:0] n2314_o;
  wire [33:0] n2316_o;
  wire [127:0] n2319_o;
  reg [33:0] n2320_q;
  wire [31:0] n2321_o;
  wire [31:0] n2322_o;
  wire [31:0] n2323_o;
  wire [31:0] n2324_o;
  wire [1:0] n2325_o;
  reg [31:0] n2326_o;
  assign bus_rsp_o_data = n2125_o; //(module output)
  assign bus_rsp_o_ack = n2126_o; //(module output)
  assign bus_rsp_o_err = n2127_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:50:5  */
  assign n2123_o = {bus_req_i_fence, bus_req_i_rvso, bus_req_i_priv, bus_req_i_src, bus_req_i_rw, bus_req_i_stb, bus_req_i_ben, bus_req_i_data, bus_req_i_addr};
  assign n2125_o = n2320_q[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:143:3  */
  assign n2126_o = n2320_q[32]; // extract
  assign n2127_o = n2320_q[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:106:10  */
  assign sysinfo = n2319_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:122:25  */
  assign n2138_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:123:25  */
  assign n2142_o = 1'b1 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:124:25  */
  assign n2146_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:125:25  */
  assign n2150_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:126:25  */
  assign n2154_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:127:25  */
  assign n2158_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:128:25  */
  assign n2162_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:129:25  */
  assign n2166_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:130:25  */
  assign n2170_o = 1'b1 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:131:25  */
  assign n2174_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:132:25  */
  assign n2178_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:136:25  */
  assign n2185_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:137:25  */
  assign n2189_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:138:25  */
  assign n2193_o = 1'b1 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:139:25  */
  assign n2197_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:140:25  */
  assign n2201_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:141:25  */
  assign n2205_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:142:25  */
  assign n2209_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:143:25  */
  assign n2213_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:144:25  */
  assign n2217_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:145:25  */
  assign n2221_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:146:25  */
  assign n2225_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:147:25  */
  assign n2229_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:148:25  */
  assign n2233_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:149:25  */
  assign n2237_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:150:25  */
  assign n2241_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:151:25  */
  assign n2245_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:152:25  */
  assign n2249_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:153:25  */
  assign n2253_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:156:98  */
  assign n2258_o = 1'b0 ? 4'b0110 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:157:98  */
  assign n2263_o = 1'b0 ? 4'b0010 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:159:98  */
  assign n2268_o = 1'b0 ? 4'b0110 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:160:98  */
  assign n2273_o = 1'b0 ? 4'b0010 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:162:101  */
  assign n2277_o = 1'b0 ? 4'b1000 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:163:101  */
  assign n2281_o = 1'b0 ? 4'b0011 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:165:102  */
  assign n2285_o = 1'b1 ? 4'b0101 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:166:102  */
  assign n2289_o = 1'b1 ? 4'b0101 : 4'b0000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:173:16  */
  assign n2292_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:181:21  */
  assign n2300_o = n2123_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:181:47  */
  assign n2301_o = n2123_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:181:50  */
  assign n2302_o = ~n2301_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:181:32  */
  assign n2303_o = n2302_o & n2300_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:183:69  */
  assign n2305_o = n2123_o[3:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:183:35  */
  assign n2308_o = 2'b11 - n2305_o;
  assign n2311_o = {1'b1, n2326_o};
  assign n2312_o = {1'b0, 32'b00000000000000000000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:181:7  */
  assign n2313_o = n2303_o ? n2311_o : n2312_o;
  assign n2314_o = {1'b0, n2313_o};
  assign n2316_o = {1'b0, 1'b0, 32'b00000000000000000000000000000000};
  assign n2319_o = {32'b00000000000000000000000000000000, 8'b00000010, 8'b00000000, 8'b00001101, 8'b00001110, n2253_o, n2249_o, n2245_o, n2241_o, n2237_o, n2233_o, n2229_o, n2225_o, n2221_o, n2217_o, n2213_o, n2209_o, n2205_o, n2201_o, n2197_o, n2193_o, n2189_o, n2185_o, 1'b0, 1'b0, 1'b0, n2178_o, n2174_o, n2170_o, n2166_o, n2162_o, n2158_o, n2154_o, n2150_o, n2146_o, n2142_o, n2138_o, n2289_o, n2285_o, n2281_o, n2277_o, n2273_o, n2268_o, n2263_o, n2258_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:177:5  */
  always @(posedge clk_i or posedge n2292_o)
    if (n2292_o)
      n2320_q <= n2316_o;
    else
      n2320_q <= n2314_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:92:5  */
  assign n2321_o = sysinfo[31:0]; // extract
  assign n2322_o = sysinfo[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:183:35  */
  assign n2323_o = sysinfo[95:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:171:3  */
  assign n2324_o = sysinfo[127:96]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:183:34  */
  assign n2325_o = n2308_o[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_sysinfo.vhd:183:34  */
  always @*
    case (n2325_o)
      2'b00: n2326_o = n2321_o;
      2'b01: n2326_o = n2322_o;
      2'b10: n2326_o = n2323_o;
      2'b11: n2326_o = n2324_o;
    endcase
endmodule

module neorv32_mtime
  (input  clk_i,
   input  rstn_i,
   input  [31:0] bus_req_i_addr,
   input  [31:0] bus_req_i_data,
   input  [3:0] bus_req_i_ben,
   input  bus_req_i_stb,
   input  bus_req_i_rw,
   input  bus_req_i_src,
   input  bus_req_i_priv,
   input  bus_req_i_rvso,
   input  bus_req_i_fence,
   output [31:0] bus_rsp_o_data,
   output bus_rsp_o_ack,
   output bus_rsp_o_err,
   output [63:0] time_o,
   output irq_o);
  wire [73:0] n1989_o;
  wire [31:0] n1991_o;
  wire n1992_o;
  wire n1993_o;
  wire [1:0] mtime_we;
  wire [31:0] mtimecmp_lo;
  wire [31:0] mtimecmp_hi;
  wire [31:0] mtime_lo;
  wire [32:0] mtime_lo_nxt;
  wire mtime_lo_cry;
  wire [31:0] mtime_hi;
  wire cmp_lo_ge;
  wire cmp_lo_ge_ff;
  wire cmp_hi_eq;
  wire cmp_hi_gt;
  wire n1997_o;
  wire n2002_o;
  wire n2003_o;
  wire n2004_o;
  wire n2005_o;
  wire n2006_o;
  wire n2007_o;
  wire n2008_o;
  wire [31:0] n2009_o;
  wire [31:0] n2010_o;
  wire [31:0] n2012_o;
  wire n2013_o;
  wire n2015_o;
  wire n2016_o;
  wire n2017_o;
  wire n2018_o;
  wire n2019_o;
  wire n2020_o;
  wire n2021_o;
  wire n2022_o;
  wire n2023_o;
  wire n2024_o;
  wire n2025_o;
  wire n2026_o;
  wire n2027_o;
  wire n2028_o;
  wire n2029_o;
  wire n2030_o;
  wire n2031_o;
  wire n2032_o;
  wire [31:0] n2033_o;
  wire [31:0] n2034_o;
  wire [31:0] n2035_o;
  wire n2036_o;
  wire n2037_o;
  wire [31:0] n2038_o;
  wire [31:0] n2039_o;
  wire [31:0] n2040_o;
  wire [31:0] n2041_o;
  wire n2042_o;
  wire n2045_o;
  wire n2046_o;
  wire n2047_o;
  wire n2048_o;
  wire [1:0] n2049_o;
  wire n2051_o;
  wire n2053_o;
  wire n2055_o;
  wire [2:0] n2056_o;
  reg [31:0] n2057_o;
  wire [31:0] n2058_o;
  wire [33:0] n2059_o;
  wire [1:0] n2061_o;
  wire [33:0] n2068_o;
  wire [32:0] n2084_o;
  wire [32:0] n2086_o;
  wire [63:0] n2087_o;
  wire n2089_o;
  wire n2091_o;
  wire n2092_o;
  wire n2101_o;
  wire n2102_o;
  wire n2105_o;
  wire n2106_o;
  wire n2109_o;
  wire n2110_o;
  reg [1:0] n2112_q;
  wire [31:0] n2113_o;
  reg [31:0] n2114_q;
  wire [31:0] n2115_o;
  reg [31:0] n2116_q;
  reg [31:0] n2117_q;
  reg n2118_q;
  reg [31:0] n2119_q;
  reg n2120_q;
  reg [33:0] n2121_q;
  reg n2122_q;
  assign bus_rsp_o_data = n1991_o; //(module output)
  assign bus_rsp_o_ack = n1992_o; //(module output)
  assign bus_rsp_o_err = n1993_o; //(module output)
  assign time_o = n2087_o; //(module output)
  assign irq_o = n2122_q; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:481:5  */
  assign n1989_o = {bus_req_i_fence, bus_req_i_rvso, bus_req_i_priv, bus_req_i_src, bus_req_i_rw, bus_req_i_stb, bus_req_i_ben, bus_req_i_data, bus_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:479:5  */
  assign n1991_o = n2121_q[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:478:5  */
  assign n1992_o = n2121_q[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:477:5  */
  assign n1993_o = n2121_q[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:58:10  */
  assign mtime_we = n2112_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:61:10  */
  assign mtimecmp_lo = n2114_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:62:10  */
  assign mtimecmp_hi = n2116_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:63:10  */
  assign mtime_lo = n2117_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:64:10  */
  assign mtime_lo_nxt = n2086_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:65:10  */
  assign mtime_lo_cry = n2118_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:66:10  */
  assign mtime_hi = n2119_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:69:10  */
  assign cmp_lo_ge = n2102_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:69:21  */
  assign cmp_lo_ge_ff = n2120_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:69:35  */
  assign cmp_hi_eq = n2106_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:69:46  */
  assign cmp_hi_gt = n2110_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:77:16  */
  assign n1997_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:90:21  */
  assign n2002_o = n1989_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:90:47  */
  assign n2003_o = n1989_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:90:32  */
  assign n2004_o = n2003_o & n2002_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:90:76  */
  assign n2005_o = n1989_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:90:57  */
  assign n2006_o = n2005_o & n2004_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:91:27  */
  assign n2007_o = n1989_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:91:31  */
  assign n2008_o = ~n2007_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:92:36  */
  assign n2009_o = n1989_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:94:36  */
  assign n2010_o = n1989_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:91:9  */
  assign n2012_o = n2008_o ? mtimecmp_hi : n2010_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:90:7  */
  assign n2013_o = n2008_o & n2006_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:32  */
  assign n2015_o = n1989_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:50  */
  assign n2016_o = n1989_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:36  */
  assign n2017_o = n2015_o & n2016_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:76  */
  assign n2018_o = n1989_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:58  */
  assign n2019_o = ~n2018_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:53  */
  assign n2020_o = n2017_o & n2019_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:104  */
  assign n2021_o = n1989_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:86  */
  assign n2022_o = ~n2021_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:99:81  */
  assign n2023_o = n2020_o & n2022_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:100:32  */
  assign n2024_o = n1989_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:100:50  */
  assign n2025_o = n1989_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:100:36  */
  assign n2026_o = n2024_o & n2025_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:100:76  */
  assign n2027_o = n1989_o[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:100:58  */
  assign n2028_o = ~n2027_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:100:53  */
  assign n2029_o = n2026_o & n2028_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:100:104  */
  assign n2030_o = n1989_o[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:100:81  */
  assign n2031_o = n2029_o & n2030_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:103:19  */
  assign n2032_o = mtime_we[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:104:31  */
  assign n2033_o = n1989_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:106:33  */
  assign n2034_o = mtime_lo_nxt[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:103:7  */
  assign n2035_o = n2032_o ? n2033_o : n2034_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:110:38  */
  assign n2036_o = mtime_lo_nxt[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:113:19  */
  assign n2037_o = mtime_we[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:114:31  */
  assign n2038_o = n1989_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:116:58  */
  assign n2039_o = {31'b0, mtime_lo_cry};  //  uext
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:116:58  */
  assign n2040_o = mtime_hi + n2039_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:113:7  */
  assign n2041_o = n2037_o ? n2038_o : n2040_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:120:35  */
  assign n2042_o = n1989_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:123:21  */
  assign n2045_o = n1989_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:123:47  */
  assign n2046_o = n1989_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:123:50  */
  assign n2047_o = ~n2046_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:123:32  */
  assign n2048_o = n2047_o & n2045_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:124:28  */
  assign n2049_o = n1989_o[3:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:125:11  */
  assign n2051_o = n2049_o == 2'b00;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:126:11  */
  assign n2053_o = n2049_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:127:11  */
  assign n2055_o = n2049_o == 2'b10;
  assign n2056_o = {n2055_o, n2053_o, n2051_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:124:9  */
  always @*
    case (n2056_o)
      3'b100: n2057_o = mtimecmp_lo;
      3'b010: n2057_o = mtime_hi;
      3'b001: n2057_o = mtime_lo;
      default: n2057_o = mtimecmp_hi;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:123:7  */
  assign n2058_o = n2048_o ? n2057_o : 32'b00000000000000000000000000000000;
  assign n2059_o = {1'b0, n2042_o, n2058_o};
  assign n2061_o = {n2031_o, n2023_o};
  assign n2068_o = {1'b0, 1'b0, 32'b00000000000000000000000000000000};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:135:50  */
  assign n2084_o = {1'b0, mtime_lo};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:135:62  */
  assign n2086_o = n2084_o + 33'b000000000000000000000000000000001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:138:22  */
  assign n2087_o = {mtime_hi, mtime_lo};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:145:16  */
  assign n2089_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:150:47  */
  assign n2091_o = cmp_hi_eq & cmp_lo_ge_ff;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:150:33  */
  assign n2092_o = cmp_hi_gt | n2091_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:155:45  */
  assign n2101_o = $unsigned(mtime_lo) >= $unsigned(mtimecmp_lo);
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:155:20  */
  assign n2102_o = n2101_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:156:45  */
  assign n2105_o = mtime_hi == mtimecmp_hi;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:156:20  */
  assign n2106_o = n2105_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:157:45  */
  assign n2109_o = $unsigned(mtime_hi) > $unsigned(mtimecmp_hi);
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:157:20  */
  assign n2110_o = n2109_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  always @(posedge clk_i or posedge n1997_o)
    if (n1997_o)
      n2112_q <= 2'b00;
    else
      n2112_q <= n2061_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  assign n2113_o = n2013_o ? n2009_o : mtimecmp_lo;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  always @(posedge clk_i or posedge n1997_o)
    if (n1997_o)
      n2114_q <= 32'b00000000000000000000000000000000;
    else
      n2114_q <= n2113_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  assign n2115_o = n2006_o ? n2012_o : mtimecmp_hi;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  always @(posedge clk_i or posedge n1997_o)
    if (n1997_o)
      n2116_q <= 32'b00000000000000000000000000000000;
    else
      n2116_q <= n2115_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  always @(posedge clk_i or posedge n1997_o)
    if (n1997_o)
      n2117_q <= 32'b00000000000000000000000000000000;
    else
      n2117_q <= n2035_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  always @(posedge clk_i or posedge n1997_o)
    if (n1997_o)
      n2118_q <= 1'b0;
    else
      n2118_q <= n2036_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  always @(posedge clk_i or posedge n1997_o)
    if (n1997_o)
      n2119_q <= 32'b00000000000000000000000000000000;
    else
      n2119_q <= n2041_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:148:5  */
  always @(posedge clk_i or posedge n2089_o)
    if (n2089_o)
      n2120_q <= 1'b0;
    else
      n2120_q <= cmp_lo_ge;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:88:5  */
  always @(posedge clk_i or posedge n1997_o)
    if (n1997_o)
      n2121_q <= n2068_o;
    else
      n2121_q <= n2059_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_mtime.vhd:148:5  */
  always @(posedge clk_i or posedge n2089_o)
    if (n2089_o)
      n2122_q <= 1'b0;
    else
      n2122_q <= n2092_o;
endmodule

module neorv32_bus_io_switch_256_84bc3e102e5c7d00d4cf85e98418cab7f8480bb6
  (input  [31:0] main_req_i_addr,
   input  [31:0] main_req_i_data,
   input  [3:0] main_req_i_ben,
   input  main_req_i_stb,
   input  main_req_i_rw,
   input  main_req_i_src,
   input  main_req_i_priv,
   input  main_req_i_rvso,
   input  main_req_i_fence,
   input  [31:0] dev_00_rsp_i_data,
   input  dev_00_rsp_i_ack,
   input  dev_00_rsp_i_err,
   input  [31:0] dev_01_rsp_i_data,
   input  dev_01_rsp_i_ack,
   input  dev_01_rsp_i_err,
   input  [31:0] dev_02_rsp_i_data,
   input  dev_02_rsp_i_ack,
   input  dev_02_rsp_i_err,
   input  [31:0] dev_03_rsp_i_data,
   input  dev_03_rsp_i_ack,
   input  dev_03_rsp_i_err,
   input  [31:0] dev_04_rsp_i_data,
   input  dev_04_rsp_i_ack,
   input  dev_04_rsp_i_err,
   input  [31:0] dev_05_rsp_i_data,
   input  dev_05_rsp_i_ack,
   input  dev_05_rsp_i_err,
   input  [31:0] dev_06_rsp_i_data,
   input  dev_06_rsp_i_ack,
   input  dev_06_rsp_i_err,
   input  [31:0] dev_07_rsp_i_data,
   input  dev_07_rsp_i_ack,
   input  dev_07_rsp_i_err,
   input  [31:0] dev_08_rsp_i_data,
   input  dev_08_rsp_i_ack,
   input  dev_08_rsp_i_err,
   input  [31:0] dev_09_rsp_i_data,
   input  dev_09_rsp_i_ack,
   input  dev_09_rsp_i_err,
   input  [31:0] dev_10_rsp_i_data,
   input  dev_10_rsp_i_ack,
   input  dev_10_rsp_i_err,
   input  [31:0] dev_11_rsp_i_data,
   input  dev_11_rsp_i_ack,
   input  dev_11_rsp_i_err,
   input  [31:0] dev_12_rsp_i_data,
   input  dev_12_rsp_i_ack,
   input  dev_12_rsp_i_err,
   input  [31:0] dev_13_rsp_i_data,
   input  dev_13_rsp_i_ack,
   input  dev_13_rsp_i_err,
   input  [31:0] dev_14_rsp_i_data,
   input  dev_14_rsp_i_ack,
   input  dev_14_rsp_i_err,
   input  [31:0] dev_15_rsp_i_data,
   input  dev_15_rsp_i_ack,
   input  dev_15_rsp_i_err,
   input  [31:0] dev_16_rsp_i_data,
   input  dev_16_rsp_i_ack,
   input  dev_16_rsp_i_err,
   input  [31:0] dev_17_rsp_i_data,
   input  dev_17_rsp_i_ack,
   input  dev_17_rsp_i_err,
   input  [31:0] dev_18_rsp_i_data,
   input  dev_18_rsp_i_ack,
   input  dev_18_rsp_i_err,
   input  [31:0] dev_19_rsp_i_data,
   input  dev_19_rsp_i_ack,
   input  dev_19_rsp_i_err,
   input  [31:0] dev_20_rsp_i_data,
   input  dev_20_rsp_i_ack,
   input  dev_20_rsp_i_err,
   output [31:0] main_rsp_o_data,
   output main_rsp_o_ack,
   output main_rsp_o_err,
   output [31:0] dev_00_req_o_addr,
   output [31:0] dev_00_req_o_data,
   output [3:0] dev_00_req_o_ben,
   output dev_00_req_o_stb,
   output dev_00_req_o_rw,
   output dev_00_req_o_src,
   output dev_00_req_o_priv,
   output dev_00_req_o_rvso,
   output dev_00_req_o_fence,
   output [31:0] dev_01_req_o_addr,
   output [31:0] dev_01_req_o_data,
   output [3:0] dev_01_req_o_ben,
   output dev_01_req_o_stb,
   output dev_01_req_o_rw,
   output dev_01_req_o_src,
   output dev_01_req_o_priv,
   output dev_01_req_o_rvso,
   output dev_01_req_o_fence,
   output [31:0] dev_02_req_o_addr,
   output [31:0] dev_02_req_o_data,
   output [3:0] dev_02_req_o_ben,
   output dev_02_req_o_stb,
   output dev_02_req_o_rw,
   output dev_02_req_o_src,
   output dev_02_req_o_priv,
   output dev_02_req_o_rvso,
   output dev_02_req_o_fence,
   output [31:0] dev_03_req_o_addr,
   output [31:0] dev_03_req_o_data,
   output [3:0] dev_03_req_o_ben,
   output dev_03_req_o_stb,
   output dev_03_req_o_rw,
   output dev_03_req_o_src,
   output dev_03_req_o_priv,
   output dev_03_req_o_rvso,
   output dev_03_req_o_fence,
   output [31:0] dev_04_req_o_addr,
   output [31:0] dev_04_req_o_data,
   output [3:0] dev_04_req_o_ben,
   output dev_04_req_o_stb,
   output dev_04_req_o_rw,
   output dev_04_req_o_src,
   output dev_04_req_o_priv,
   output dev_04_req_o_rvso,
   output dev_04_req_o_fence,
   output [31:0] dev_05_req_o_addr,
   output [31:0] dev_05_req_o_data,
   output [3:0] dev_05_req_o_ben,
   output dev_05_req_o_stb,
   output dev_05_req_o_rw,
   output dev_05_req_o_src,
   output dev_05_req_o_priv,
   output dev_05_req_o_rvso,
   output dev_05_req_o_fence,
   output [31:0] dev_06_req_o_addr,
   output [31:0] dev_06_req_o_data,
   output [3:0] dev_06_req_o_ben,
   output dev_06_req_o_stb,
   output dev_06_req_o_rw,
   output dev_06_req_o_src,
   output dev_06_req_o_priv,
   output dev_06_req_o_rvso,
   output dev_06_req_o_fence,
   output [31:0] dev_07_req_o_addr,
   output [31:0] dev_07_req_o_data,
   output [3:0] dev_07_req_o_ben,
   output dev_07_req_o_stb,
   output dev_07_req_o_rw,
   output dev_07_req_o_src,
   output dev_07_req_o_priv,
   output dev_07_req_o_rvso,
   output dev_07_req_o_fence,
   output [31:0] dev_08_req_o_addr,
   output [31:0] dev_08_req_o_data,
   output [3:0] dev_08_req_o_ben,
   output dev_08_req_o_stb,
   output dev_08_req_o_rw,
   output dev_08_req_o_src,
   output dev_08_req_o_priv,
   output dev_08_req_o_rvso,
   output dev_08_req_o_fence,
   output [31:0] dev_09_req_o_addr,
   output [31:0] dev_09_req_o_data,
   output [3:0] dev_09_req_o_ben,
   output dev_09_req_o_stb,
   output dev_09_req_o_rw,
   output dev_09_req_o_src,
   output dev_09_req_o_priv,
   output dev_09_req_o_rvso,
   output dev_09_req_o_fence,
   output [31:0] dev_10_req_o_addr,
   output [31:0] dev_10_req_o_data,
   output [3:0] dev_10_req_o_ben,
   output dev_10_req_o_stb,
   output dev_10_req_o_rw,
   output dev_10_req_o_src,
   output dev_10_req_o_priv,
   output dev_10_req_o_rvso,
   output dev_10_req_o_fence,
   output [31:0] dev_11_req_o_addr,
   output [31:0] dev_11_req_o_data,
   output [3:0] dev_11_req_o_ben,
   output dev_11_req_o_stb,
   output dev_11_req_o_rw,
   output dev_11_req_o_src,
   output dev_11_req_o_priv,
   output dev_11_req_o_rvso,
   output dev_11_req_o_fence,
   output [31:0] dev_12_req_o_addr,
   output [31:0] dev_12_req_o_data,
   output [3:0] dev_12_req_o_ben,
   output dev_12_req_o_stb,
   output dev_12_req_o_rw,
   output dev_12_req_o_src,
   output dev_12_req_o_priv,
   output dev_12_req_o_rvso,
   output dev_12_req_o_fence,
   output [31:0] dev_13_req_o_addr,
   output [31:0] dev_13_req_o_data,
   output [3:0] dev_13_req_o_ben,
   output dev_13_req_o_stb,
   output dev_13_req_o_rw,
   output dev_13_req_o_src,
   output dev_13_req_o_priv,
   output dev_13_req_o_rvso,
   output dev_13_req_o_fence,
   output [31:0] dev_14_req_o_addr,
   output [31:0] dev_14_req_o_data,
   output [3:0] dev_14_req_o_ben,
   output dev_14_req_o_stb,
   output dev_14_req_o_rw,
   output dev_14_req_o_src,
   output dev_14_req_o_priv,
   output dev_14_req_o_rvso,
   output dev_14_req_o_fence,
   output [31:0] dev_15_req_o_addr,
   output [31:0] dev_15_req_o_data,
   output [3:0] dev_15_req_o_ben,
   output dev_15_req_o_stb,
   output dev_15_req_o_rw,
   output dev_15_req_o_src,
   output dev_15_req_o_priv,
   output dev_15_req_o_rvso,
   output dev_15_req_o_fence,
   output [31:0] dev_16_req_o_addr,
   output [31:0] dev_16_req_o_data,
   output [3:0] dev_16_req_o_ben,
   output dev_16_req_o_stb,
   output dev_16_req_o_rw,
   output dev_16_req_o_src,
   output dev_16_req_o_priv,
   output dev_16_req_o_rvso,
   output dev_16_req_o_fence,
   output [31:0] dev_17_req_o_addr,
   output [31:0] dev_17_req_o_data,
   output [3:0] dev_17_req_o_ben,
   output dev_17_req_o_stb,
   output dev_17_req_o_rw,
   output dev_17_req_o_src,
   output dev_17_req_o_priv,
   output dev_17_req_o_rvso,
   output dev_17_req_o_fence,
   output [31:0] dev_18_req_o_addr,
   output [31:0] dev_18_req_o_data,
   output [3:0] dev_18_req_o_ben,
   output dev_18_req_o_stb,
   output dev_18_req_o_rw,
   output dev_18_req_o_src,
   output dev_18_req_o_priv,
   output dev_18_req_o_rvso,
   output dev_18_req_o_fence,
   output [31:0] dev_19_req_o_addr,
   output [31:0] dev_19_req_o_data,
   output [3:0] dev_19_req_o_ben,
   output dev_19_req_o_stb,
   output dev_19_req_o_rw,
   output dev_19_req_o_src,
   output dev_19_req_o_priv,
   output dev_19_req_o_rvso,
   output dev_19_req_o_fence,
   output [31:0] dev_20_req_o_addr,
   output [31:0] dev_20_req_o_data,
   output [3:0] dev_20_req_o_ben,
   output dev_20_req_o_stb,
   output dev_20_req_o_rw,
   output dev_20_req_o_src,
   output dev_20_req_o_priv,
   output dev_20_req_o_rvso,
   output dev_20_req_o_fence);
  wire [73:0] n1671_o;
  wire [31:0] n1673_o;
  wire n1674_o;
  wire n1675_o;
  wire [31:0] n1677_o;
  wire [31:0] n1678_o;
  wire [3:0] n1679_o;
  wire n1680_o;
  wire n1681_o;
  wire n1682_o;
  wire n1683_o;
  wire n1684_o;
  wire n1685_o;
  wire [33:0] n1686_o;
  wire [31:0] n1688_o;
  wire [31:0] n1689_o;
  wire [3:0] n1690_o;
  wire n1691_o;
  wire n1692_o;
  wire n1693_o;
  wire n1694_o;
  wire n1695_o;
  wire n1696_o;
  wire [33:0] n1697_o;
  wire [31:0] n1699_o;
  wire [31:0] n1700_o;
  wire [3:0] n1701_o;
  wire n1702_o;
  wire n1703_o;
  wire n1704_o;
  wire n1705_o;
  wire n1706_o;
  wire n1707_o;
  wire [33:0] n1708_o;
  wire [31:0] n1710_o;
  wire [31:0] n1711_o;
  wire [3:0] n1712_o;
  wire n1713_o;
  wire n1714_o;
  wire n1715_o;
  wire n1716_o;
  wire n1717_o;
  wire n1718_o;
  wire [33:0] n1719_o;
  wire [31:0] n1721_o;
  wire [31:0] n1722_o;
  wire [3:0] n1723_o;
  wire n1724_o;
  wire n1725_o;
  wire n1726_o;
  wire n1727_o;
  wire n1728_o;
  wire n1729_o;
  wire [33:0] n1730_o;
  wire [31:0] n1732_o;
  wire [31:0] n1733_o;
  wire [3:0] n1734_o;
  wire n1735_o;
  wire n1736_o;
  wire n1737_o;
  wire n1738_o;
  wire n1739_o;
  wire n1740_o;
  wire [33:0] n1741_o;
  wire [31:0] n1743_o;
  wire [31:0] n1744_o;
  wire [3:0] n1745_o;
  wire n1746_o;
  wire n1747_o;
  wire n1748_o;
  wire n1749_o;
  wire n1750_o;
  wire n1751_o;
  wire [33:0] n1752_o;
  wire [31:0] n1754_o;
  wire [31:0] n1755_o;
  wire [3:0] n1756_o;
  wire n1757_o;
  wire n1758_o;
  wire n1759_o;
  wire n1760_o;
  wire n1761_o;
  wire n1762_o;
  wire [33:0] n1763_o;
  wire [31:0] n1765_o;
  wire [31:0] n1766_o;
  wire [3:0] n1767_o;
  wire n1768_o;
  wire n1769_o;
  wire n1770_o;
  wire n1771_o;
  wire n1772_o;
  wire n1773_o;
  wire [33:0] n1774_o;
  wire [31:0] n1776_o;
  wire [31:0] n1777_o;
  wire [3:0] n1778_o;
  wire n1779_o;
  wire n1780_o;
  wire n1781_o;
  wire n1782_o;
  wire n1783_o;
  wire n1784_o;
  wire [33:0] n1785_o;
  wire [31:0] n1787_o;
  wire [31:0] n1788_o;
  wire [3:0] n1789_o;
  wire n1790_o;
  wire n1791_o;
  wire n1792_o;
  wire n1793_o;
  wire n1794_o;
  wire n1795_o;
  wire [33:0] n1796_o;
  wire [31:0] n1798_o;
  wire [31:0] n1799_o;
  wire [3:0] n1800_o;
  wire n1801_o;
  wire n1802_o;
  wire n1803_o;
  wire n1804_o;
  wire n1805_o;
  wire n1806_o;
  wire [33:0] n1807_o;
  wire [31:0] n1809_o;
  wire [31:0] n1810_o;
  wire [3:0] n1811_o;
  wire n1812_o;
  wire n1813_o;
  wire n1814_o;
  wire n1815_o;
  wire n1816_o;
  wire n1817_o;
  wire [33:0] n1818_o;
  wire [31:0] n1820_o;
  wire [31:0] n1821_o;
  wire [3:0] n1822_o;
  wire n1823_o;
  wire n1824_o;
  wire n1825_o;
  wire n1826_o;
  wire n1827_o;
  wire n1828_o;
  wire [33:0] n1829_o;
  wire [31:0] n1831_o;
  wire [31:0] n1832_o;
  wire [3:0] n1833_o;
  wire n1834_o;
  wire n1835_o;
  wire n1836_o;
  wire n1837_o;
  wire n1838_o;
  wire n1839_o;
  wire [33:0] n1840_o;
  wire [31:0] n1842_o;
  wire [31:0] n1843_o;
  wire [3:0] n1844_o;
  wire n1845_o;
  wire n1846_o;
  wire n1847_o;
  wire n1848_o;
  wire n1849_o;
  wire n1850_o;
  wire [33:0] n1851_o;
  wire [31:0] n1853_o;
  wire [31:0] n1854_o;
  wire [3:0] n1855_o;
  wire n1856_o;
  wire n1857_o;
  wire n1858_o;
  wire n1859_o;
  wire n1860_o;
  wire n1861_o;
  wire [33:0] n1862_o;
  wire [31:0] n1864_o;
  wire [31:0] n1865_o;
  wire [3:0] n1866_o;
  wire n1867_o;
  wire n1868_o;
  wire n1869_o;
  wire n1870_o;
  wire n1871_o;
  wire n1872_o;
  wire [33:0] n1873_o;
  wire [31:0] n1875_o;
  wire [31:0] n1876_o;
  wire [3:0] n1877_o;
  wire n1878_o;
  wire n1879_o;
  wire n1880_o;
  wire n1881_o;
  wire n1882_o;
  wire n1883_o;
  wire [33:0] n1884_o;
  wire [31:0] n1886_o;
  wire [31:0] n1887_o;
  wire [3:0] n1888_o;
  wire n1889_o;
  wire n1890_o;
  wire n1891_o;
  wire n1892_o;
  wire n1893_o;
  wire n1894_o;
  wire [33:0] n1895_o;
  wire [31:0] n1897_o;
  wire [31:0] n1898_o;
  wire [3:0] n1899_o;
  wire n1900_o;
  wire n1901_o;
  wire n1902_o;
  wire n1903_o;
  wire n1904_o;
  wire n1905_o;
  wire [33:0] n1906_o;
  wire [1553:0] dev_req;
  wire [713:0] dev_rsp;
  wire [73:0] n1907_o;
  wire [73:0] n1908_o;
  wire [73:0] n1909_o;
  wire [73:0] n1910_o;
  wire [73:0] n1911_o;
  wire [73:0] n1912_o;
  wire [73:0] n1913_o;
  wire [73:0] n1914_o;
  wire [73:0] n1915_o;
  wire [73:0] n1916_o;
  wire [73:0] n1917_o;
  wire [73:0] n1918_o;
  wire [73:0] n1919_o;
  wire [73:0] n1920_o;
  wire [73:0] n1921_o;
  wire [73:0] n1922_o;
  wire [73:0] n1923_o;
  wire [73:0] n1924_o;
  wire [73:0] n1925_o;
  wire [73:0] n1926_o;
  wire [73:0] n1927_o;
  wire [4:0] n1930_o;
  wire n1932_o;
  wire n1933_o;
  wire n1935_o;
  wire [4:0] n1936_o;
  wire [67:0] n1937_o;
  wire [4:0] n1940_o;
  wire n1942_o;
  wire n1943_o;
  wire n1945_o;
  wire [4:0] n1946_o;
  wire [67:0] n1947_o;
  localparam [33:0] n1951_o = 34'b0000000000000000000000000000000000;
  wire [31:0] n1952_o;
  wire [31:0] n1954_o;
  wire [31:0] n1955_o;
  localparam [33:0] n1956_o = 34'b0000000000000000000000000000000000;
  wire [1:0] n1957_o;
  wire [33:0] n1958_o;
  wire n1959_o;
  wire n1961_o;
  wire n1962_o;
  wire n1963_o;
  wire [33:0] n1964_o;
  wire n1965_o;
  wire n1967_o;
  wire n1968_o;
  wire [33:0] n1969_o;
  wire [31:0] n1970_o;
  wire [31:0] n1972_o;
  wire [31:0] n1973_o;
  wire [33:0] n1974_o;
  wire n1975_o;
  wire n1977_o;
  wire n1978_o;
  wire [33:0] n1979_o;
  wire n1980_o;
  wire n1982_o;
  wire n1983_o;
  wire [33:0] n1984_o;
  wire [1553:0] n1987_o;
  wire [713:0] n1988_o;
  assign main_rsp_o_data = n1673_o; //(module output)
  assign main_rsp_o_ack = n1674_o; //(module output)
  assign main_rsp_o_err = n1675_o; //(module output)
  assign dev_00_req_o_addr = n1677_o; //(module output)
  assign dev_00_req_o_data = n1678_o; //(module output)
  assign dev_00_req_o_ben = n1679_o; //(module output)
  assign dev_00_req_o_stb = n1680_o; //(module output)
  assign dev_00_req_o_rw = n1681_o; //(module output)
  assign dev_00_req_o_src = n1682_o; //(module output)
  assign dev_00_req_o_priv = n1683_o; //(module output)
  assign dev_00_req_o_rvso = n1684_o; //(module output)
  assign dev_00_req_o_fence = n1685_o; //(module output)
  assign dev_01_req_o_addr = n1688_o; //(module output)
  assign dev_01_req_o_data = n1689_o; //(module output)
  assign dev_01_req_o_ben = n1690_o; //(module output)
  assign dev_01_req_o_stb = n1691_o; //(module output)
  assign dev_01_req_o_rw = n1692_o; //(module output)
  assign dev_01_req_o_src = n1693_o; //(module output)
  assign dev_01_req_o_priv = n1694_o; //(module output)
  assign dev_01_req_o_rvso = n1695_o; //(module output)
  assign dev_01_req_o_fence = n1696_o; //(module output)
  assign dev_02_req_o_addr = n1699_o; //(module output)
  assign dev_02_req_o_data = n1700_o; //(module output)
  assign dev_02_req_o_ben = n1701_o; //(module output)
  assign dev_02_req_o_stb = n1702_o; //(module output)
  assign dev_02_req_o_rw = n1703_o; //(module output)
  assign dev_02_req_o_src = n1704_o; //(module output)
  assign dev_02_req_o_priv = n1705_o; //(module output)
  assign dev_02_req_o_rvso = n1706_o; //(module output)
  assign dev_02_req_o_fence = n1707_o; //(module output)
  assign dev_03_req_o_addr = n1710_o; //(module output)
  assign dev_03_req_o_data = n1711_o; //(module output)
  assign dev_03_req_o_ben = n1712_o; //(module output)
  assign dev_03_req_o_stb = n1713_o; //(module output)
  assign dev_03_req_o_rw = n1714_o; //(module output)
  assign dev_03_req_o_src = n1715_o; //(module output)
  assign dev_03_req_o_priv = n1716_o; //(module output)
  assign dev_03_req_o_rvso = n1717_o; //(module output)
  assign dev_03_req_o_fence = n1718_o; //(module output)
  assign dev_04_req_o_addr = n1721_o; //(module output)
  assign dev_04_req_o_data = n1722_o; //(module output)
  assign dev_04_req_o_ben = n1723_o; //(module output)
  assign dev_04_req_o_stb = n1724_o; //(module output)
  assign dev_04_req_o_rw = n1725_o; //(module output)
  assign dev_04_req_o_src = n1726_o; //(module output)
  assign dev_04_req_o_priv = n1727_o; //(module output)
  assign dev_04_req_o_rvso = n1728_o; //(module output)
  assign dev_04_req_o_fence = n1729_o; //(module output)
  assign dev_05_req_o_addr = n1732_o; //(module output)
  assign dev_05_req_o_data = n1733_o; //(module output)
  assign dev_05_req_o_ben = n1734_o; //(module output)
  assign dev_05_req_o_stb = n1735_o; //(module output)
  assign dev_05_req_o_rw = n1736_o; //(module output)
  assign dev_05_req_o_src = n1737_o; //(module output)
  assign dev_05_req_o_priv = n1738_o; //(module output)
  assign dev_05_req_o_rvso = n1739_o; //(module output)
  assign dev_05_req_o_fence = n1740_o; //(module output)
  assign dev_06_req_o_addr = n1743_o; //(module output)
  assign dev_06_req_o_data = n1744_o; //(module output)
  assign dev_06_req_o_ben = n1745_o; //(module output)
  assign dev_06_req_o_stb = n1746_o; //(module output)
  assign dev_06_req_o_rw = n1747_o; //(module output)
  assign dev_06_req_o_src = n1748_o; //(module output)
  assign dev_06_req_o_priv = n1749_o; //(module output)
  assign dev_06_req_o_rvso = n1750_o; //(module output)
  assign dev_06_req_o_fence = n1751_o; //(module output)
  assign dev_07_req_o_addr = n1754_o; //(module output)
  assign dev_07_req_o_data = n1755_o; //(module output)
  assign dev_07_req_o_ben = n1756_o; //(module output)
  assign dev_07_req_o_stb = n1757_o; //(module output)
  assign dev_07_req_o_rw = n1758_o; //(module output)
  assign dev_07_req_o_src = n1759_o; //(module output)
  assign dev_07_req_o_priv = n1760_o; //(module output)
  assign dev_07_req_o_rvso = n1761_o; //(module output)
  assign dev_07_req_o_fence = n1762_o; //(module output)
  assign dev_08_req_o_addr = n1765_o; //(module output)
  assign dev_08_req_o_data = n1766_o; //(module output)
  assign dev_08_req_o_ben = n1767_o; //(module output)
  assign dev_08_req_o_stb = n1768_o; //(module output)
  assign dev_08_req_o_rw = n1769_o; //(module output)
  assign dev_08_req_o_src = n1770_o; //(module output)
  assign dev_08_req_o_priv = n1771_o; //(module output)
  assign dev_08_req_o_rvso = n1772_o; //(module output)
  assign dev_08_req_o_fence = n1773_o; //(module output)
  assign dev_09_req_o_addr = n1776_o; //(module output)
  assign dev_09_req_o_data = n1777_o; //(module output)
  assign dev_09_req_o_ben = n1778_o; //(module output)
  assign dev_09_req_o_stb = n1779_o; //(module output)
  assign dev_09_req_o_rw = n1780_o; //(module output)
  assign dev_09_req_o_src = n1781_o; //(module output)
  assign dev_09_req_o_priv = n1782_o; //(module output)
  assign dev_09_req_o_rvso = n1783_o; //(module output)
  assign dev_09_req_o_fence = n1784_o; //(module output)
  assign dev_10_req_o_addr = n1787_o; //(module output)
  assign dev_10_req_o_data = n1788_o; //(module output)
  assign dev_10_req_o_ben = n1789_o; //(module output)
  assign dev_10_req_o_stb = n1790_o; //(module output)
  assign dev_10_req_o_rw = n1791_o; //(module output)
  assign dev_10_req_o_src = n1792_o; //(module output)
  assign dev_10_req_o_priv = n1793_o; //(module output)
  assign dev_10_req_o_rvso = n1794_o; //(module output)
  assign dev_10_req_o_fence = n1795_o; //(module output)
  assign dev_11_req_o_addr = n1798_o; //(module output)
  assign dev_11_req_o_data = n1799_o; //(module output)
  assign dev_11_req_o_ben = n1800_o; //(module output)
  assign dev_11_req_o_stb = n1801_o; //(module output)
  assign dev_11_req_o_rw = n1802_o; //(module output)
  assign dev_11_req_o_src = n1803_o; //(module output)
  assign dev_11_req_o_priv = n1804_o; //(module output)
  assign dev_11_req_o_rvso = n1805_o; //(module output)
  assign dev_11_req_o_fence = n1806_o; //(module output)
  assign dev_12_req_o_addr = n1809_o; //(module output)
  assign dev_12_req_o_data = n1810_o; //(module output)
  assign dev_12_req_o_ben = n1811_o; //(module output)
  assign dev_12_req_o_stb = n1812_o; //(module output)
  assign dev_12_req_o_rw = n1813_o; //(module output)
  assign dev_12_req_o_src = n1814_o; //(module output)
  assign dev_12_req_o_priv = n1815_o; //(module output)
  assign dev_12_req_o_rvso = n1816_o; //(module output)
  assign dev_12_req_o_fence = n1817_o; //(module output)
  assign dev_13_req_o_addr = n1820_o; //(module output)
  assign dev_13_req_o_data = n1821_o; //(module output)
  assign dev_13_req_o_ben = n1822_o; //(module output)
  assign dev_13_req_o_stb = n1823_o; //(module output)
  assign dev_13_req_o_rw = n1824_o; //(module output)
  assign dev_13_req_o_src = n1825_o; //(module output)
  assign dev_13_req_o_priv = n1826_o; //(module output)
  assign dev_13_req_o_rvso = n1827_o; //(module output)
  assign dev_13_req_o_fence = n1828_o; //(module output)
  assign dev_14_req_o_addr = n1831_o; //(module output)
  assign dev_14_req_o_data = n1832_o; //(module output)
  assign dev_14_req_o_ben = n1833_o; //(module output)
  assign dev_14_req_o_stb = n1834_o; //(module output)
  assign dev_14_req_o_rw = n1835_o; //(module output)
  assign dev_14_req_o_src = n1836_o; //(module output)
  assign dev_14_req_o_priv = n1837_o; //(module output)
  assign dev_14_req_o_rvso = n1838_o; //(module output)
  assign dev_14_req_o_fence = n1839_o; //(module output)
  assign dev_15_req_o_addr = n1842_o; //(module output)
  assign dev_15_req_o_data = n1843_o; //(module output)
  assign dev_15_req_o_ben = n1844_o; //(module output)
  assign dev_15_req_o_stb = n1845_o; //(module output)
  assign dev_15_req_o_rw = n1846_o; //(module output)
  assign dev_15_req_o_src = n1847_o; //(module output)
  assign dev_15_req_o_priv = n1848_o; //(module output)
  assign dev_15_req_o_rvso = n1849_o; //(module output)
  assign dev_15_req_o_fence = n1850_o; //(module output)
  assign dev_16_req_o_addr = n1853_o; //(module output)
  assign dev_16_req_o_data = n1854_o; //(module output)
  assign dev_16_req_o_ben = n1855_o; //(module output)
  assign dev_16_req_o_stb = n1856_o; //(module output)
  assign dev_16_req_o_rw = n1857_o; //(module output)
  assign dev_16_req_o_src = n1858_o; //(module output)
  assign dev_16_req_o_priv = n1859_o; //(module output)
  assign dev_16_req_o_rvso = n1860_o; //(module output)
  assign dev_16_req_o_fence = n1861_o; //(module output)
  assign dev_17_req_o_addr = n1864_o; //(module output)
  assign dev_17_req_o_data = n1865_o; //(module output)
  assign dev_17_req_o_ben = n1866_o; //(module output)
  assign dev_17_req_o_stb = n1867_o; //(module output)
  assign dev_17_req_o_rw = n1868_o; //(module output)
  assign dev_17_req_o_src = n1869_o; //(module output)
  assign dev_17_req_o_priv = n1870_o; //(module output)
  assign dev_17_req_o_rvso = n1871_o; //(module output)
  assign dev_17_req_o_fence = n1872_o; //(module output)
  assign dev_18_req_o_addr = n1875_o; //(module output)
  assign dev_18_req_o_data = n1876_o; //(module output)
  assign dev_18_req_o_ben = n1877_o; //(module output)
  assign dev_18_req_o_stb = n1878_o; //(module output)
  assign dev_18_req_o_rw = n1879_o; //(module output)
  assign dev_18_req_o_src = n1880_o; //(module output)
  assign dev_18_req_o_priv = n1881_o; //(module output)
  assign dev_18_req_o_rvso = n1882_o; //(module output)
  assign dev_18_req_o_fence = n1883_o; //(module output)
  assign dev_19_req_o_addr = n1886_o; //(module output)
  assign dev_19_req_o_data = n1887_o; //(module output)
  assign dev_19_req_o_ben = n1888_o; //(module output)
  assign dev_19_req_o_stb = n1889_o; //(module output)
  assign dev_19_req_o_rw = n1890_o; //(module output)
  assign dev_19_req_o_src = n1891_o; //(module output)
  assign dev_19_req_o_priv = n1892_o; //(module output)
  assign dev_19_req_o_rvso = n1893_o; //(module output)
  assign dev_19_req_o_fence = n1894_o; //(module output)
  assign dev_20_req_o_addr = n1897_o; //(module output)
  assign dev_20_req_o_data = n1898_o; //(module output)
  assign dev_20_req_o_ben = n1899_o; //(module output)
  assign dev_20_req_o_stb = n1900_o; //(module output)
  assign dev_20_req_o_rw = n1901_o; //(module output)
  assign dev_20_req_o_src = n1902_o; //(module output)
  assign dev_20_req_o_priv = n1903_o; //(module output)
  assign dev_20_req_o_rvso = n1904_o; //(module output)
  assign dev_20_req_o_fence = n1905_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:381:18  */
  assign n1671_o = {main_req_i_fence, main_req_i_rvso, main_req_i_priv, main_req_i_src, main_req_i_rw, main_req_i_stb, main_req_i_ben, main_req_i_data, main_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:359:19  */
  assign n1673_o = n1984_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:358:19  */
  assign n1674_o = n1984_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:357:19  */
  assign n1675_o = n1984_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:355:19  */
  assign n1677_o = n1907_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:351:19  */
  assign n1678_o = n1907_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:350:19  */
  assign n1679_o = n1907_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:348:19  */
  assign n1680_o = n1907_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:343:19  */
  assign n1681_o = n1907_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  assign n1682_o = n1907_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  assign n1683_o = n1907_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  assign n1684_o = n1907_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  assign n1685_o = n1907_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  assign n1686_o = {dev_00_rsp_i_err, dev_00_rsp_i_ack, dev_00_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  assign n1688_o = n1908_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  assign n1689_o = n1908_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  assign n1690_o = n1908_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:321:17  */
  assign n1691_o = n1908_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:320:17  */
  assign n1692_o = n1908_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:313:17  */
  assign n1693_o = n1908_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:312:17  */
  assign n1694_o = n1908_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:311:17  */
  assign n1695_o = n1908_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:296:3  */
  assign n1696_o = n1908_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:296:3  */
  assign n1697_o = {dev_01_rsp_i_err, dev_01_rsp_i_ack, dev_01_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:296:3  */
  assign n1699_o = n1909_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:296:3  */
  assign n1700_o = n1909_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:288:19  */
  assign n1701_o = n1909_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:287:19  */
  assign n1702_o = n1909_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:286:19  */
  assign n1703_o = n1909_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:285:19  */
  assign n1704_o = n1909_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:284:19  */
  assign n1705_o = n1909_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:281:19  */
  assign n1706_o = n1909_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:278:19  */
  assign n1707_o = n1909_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:277:19  */
  assign n1708_o = {dev_02_rsp_i_err, dev_02_rsp_i_ack, dev_02_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1710_o = n1910_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1711_o = n1910_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1712_o = n1910_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1713_o = n1910_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1714_o = n1910_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1715_o = n1910_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1716_o = n1910_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1717_o = n1910_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  assign n1718_o = n1910_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:80:5  */
  assign n1719_o = {dev_03_rsp_i_err, dev_03_rsp_i_ack, dev_03_rsp_i_data};
  assign n1721_o = n1911_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:225:5  */
  assign n1722_o = n1911_o[63:32]; // extract
  assign n1723_o = n1911_o[67:64]; // extract
  assign n1724_o = n1911_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:210:3  */
  assign n1725_o = n1911_o[69]; // extract
  assign n1726_o = n1911_o[70]; // extract
  assign n1727_o = n1911_o[71]; // extract
  assign n1728_o = n1911_o[72]; // extract
  assign n1729_o = n1911_o[73]; // extract
  assign n1730_o = {dev_04_rsp_i_err, dev_04_rsp_i_ack, dev_04_rsp_i_data};
  assign n1732_o = n1912_o[31:0]; // extract
  assign n1733_o = n1912_o[63:32]; // extract
  assign n1734_o = n1912_o[67:64]; // extract
  assign n1735_o = n1912_o[68]; // extract
  assign n1736_o = n1912_o[69]; // extract
  assign n1737_o = n1912_o[70]; // extract
  assign n1738_o = n1912_o[71]; // extract
  assign n1739_o = n1912_o[72]; // extract
  assign n1740_o = n1912_o[73]; // extract
  assign n1741_o = {dev_05_rsp_i_err, dev_05_rsp_i_ack, dev_05_rsp_i_data};
  assign n1743_o = n1913_o[31:0]; // extract
  assign n1744_o = n1913_o[63:32]; // extract
  assign n1745_o = n1913_o[67:64]; // extract
  assign n1746_o = n1913_o[68]; // extract
  assign n1747_o = n1913_o[69]; // extract
  assign n1748_o = n1913_o[70]; // extract
  assign n1749_o = n1913_o[71]; // extract
  assign n1750_o = n1913_o[72]; // extract
  assign n1751_o = n1913_o[73]; // extract
  assign n1752_o = {dev_06_rsp_i_err, dev_06_rsp_i_ack, dev_06_rsp_i_data};
  assign n1754_o = n1914_o[31:0]; // extract
  assign n1755_o = n1914_o[63:32]; // extract
  assign n1756_o = n1914_o[67:64]; // extract
  assign n1757_o = n1914_o[68]; // extract
  assign n1758_o = n1914_o[69]; // extract
  assign n1759_o = n1914_o[70]; // extract
  assign n1760_o = n1914_o[71]; // extract
  assign n1761_o = n1914_o[72]; // extract
  assign n1762_o = n1914_o[73]; // extract
  assign n1763_o = {dev_07_rsp_i_err, dev_07_rsp_i_ack, dev_07_rsp_i_data};
  assign n1765_o = n1915_o[31:0]; // extract
  assign n1766_o = n1915_o[63:32]; // extract
  assign n1767_o = n1915_o[67:64]; // extract
  assign n1768_o = n1915_o[68]; // extract
  assign n1769_o = n1915_o[69]; // extract
  assign n1770_o = n1915_o[70]; // extract
  assign n1771_o = n1915_o[71]; // extract
  assign n1772_o = n1915_o[72]; // extract
  assign n1773_o = n1915_o[73]; // extract
  assign n1774_o = {dev_08_rsp_i_err, dev_08_rsp_i_ack, dev_08_rsp_i_data};
  assign n1776_o = n1916_o[31:0]; // extract
  assign n1777_o = n1916_o[63:32]; // extract
  assign n1778_o = n1916_o[67:64]; // extract
  assign n1779_o = n1916_o[68]; // extract
  assign n1780_o = n1916_o[69]; // extract
  assign n1781_o = n1916_o[70]; // extract
  assign n1782_o = n1916_o[71]; // extract
  assign n1783_o = n1916_o[72]; // extract
  assign n1784_o = n1916_o[73]; // extract
  assign n1785_o = {dev_09_rsp_i_err, dev_09_rsp_i_ack, dev_09_rsp_i_data};
  assign n1787_o = n1917_o[31:0]; // extract
  assign n1788_o = n1917_o[63:32]; // extract
  assign n1789_o = n1917_o[67:64]; // extract
  assign n1790_o = n1917_o[68]; // extract
  assign n1791_o = n1917_o[69]; // extract
  assign n1792_o = n1917_o[70]; // extract
  assign n1793_o = n1917_o[71]; // extract
  assign n1794_o = n1917_o[72]; // extract
  assign n1795_o = n1917_o[73]; // extract
  assign n1796_o = {dev_10_rsp_i_err, dev_10_rsp_i_ack, dev_10_rsp_i_data};
  assign n1798_o = n1918_o[31:0]; // extract
  assign n1799_o = n1918_o[63:32]; // extract
  assign n1800_o = n1918_o[67:64]; // extract
  assign n1801_o = n1918_o[68]; // extract
  assign n1802_o = n1918_o[69]; // extract
  assign n1803_o = n1918_o[70]; // extract
  assign n1804_o = n1918_o[71]; // extract
  assign n1805_o = n1918_o[72]; // extract
  assign n1806_o = n1918_o[73]; // extract
  assign n1807_o = {dev_11_rsp_i_err, dev_11_rsp_i_ack, dev_11_rsp_i_data};
  assign n1809_o = n1919_o[31:0]; // extract
  assign n1810_o = n1919_o[63:32]; // extract
  assign n1811_o = n1919_o[67:64]; // extract
  assign n1812_o = n1919_o[68]; // extract
  assign n1813_o = n1919_o[69]; // extract
  assign n1814_o = n1919_o[70]; // extract
  assign n1815_o = n1919_o[71]; // extract
  assign n1816_o = n1919_o[72]; // extract
  assign n1817_o = n1919_o[73]; // extract
  assign n1818_o = {dev_12_rsp_i_err, dev_12_rsp_i_ack, dev_12_rsp_i_data};
  assign n1820_o = n1920_o[31:0]; // extract
  assign n1821_o = n1920_o[63:32]; // extract
  assign n1822_o = n1920_o[67:64]; // extract
  assign n1823_o = n1920_o[68]; // extract
  assign n1824_o = n1920_o[69]; // extract
  assign n1825_o = n1920_o[70]; // extract
  assign n1826_o = n1920_o[71]; // extract
  assign n1827_o = n1920_o[72]; // extract
  assign n1828_o = n1920_o[73]; // extract
  assign n1829_o = {dev_13_rsp_i_err, dev_13_rsp_i_ack, dev_13_rsp_i_data};
  assign n1831_o = n1921_o[31:0]; // extract
  assign n1832_o = n1921_o[63:32]; // extract
  assign n1833_o = n1921_o[67:64]; // extract
  assign n1834_o = n1921_o[68]; // extract
  assign n1835_o = n1921_o[69]; // extract
  assign n1836_o = n1921_o[70]; // extract
  assign n1837_o = n1921_o[71]; // extract
  assign n1838_o = n1921_o[72]; // extract
  assign n1839_o = n1921_o[73]; // extract
  assign n1840_o = {dev_14_rsp_i_err, dev_14_rsp_i_ack, dev_14_rsp_i_data};
  assign n1842_o = n1922_o[31:0]; // extract
  assign n1843_o = n1922_o[63:32]; // extract
  assign n1844_o = n1922_o[67:64]; // extract
  assign n1845_o = n1922_o[68]; // extract
  assign n1846_o = n1922_o[69]; // extract
  assign n1847_o = n1922_o[70]; // extract
  assign n1848_o = n1922_o[71]; // extract
  assign n1849_o = n1922_o[72]; // extract
  assign n1850_o = n1922_o[73]; // extract
  assign n1851_o = {dev_15_rsp_i_err, dev_15_rsp_i_ack, dev_15_rsp_i_data};
  assign n1853_o = n1923_o[31:0]; // extract
  assign n1854_o = n1923_o[63:32]; // extract
  assign n1855_o = n1923_o[67:64]; // extract
  assign n1856_o = n1923_o[68]; // extract
  assign n1857_o = n1923_o[69]; // extract
  assign n1858_o = n1923_o[70]; // extract
  assign n1859_o = n1923_o[71]; // extract
  assign n1860_o = n1923_o[72]; // extract
  assign n1861_o = n1923_o[73]; // extract
  assign n1862_o = {dev_16_rsp_i_err, dev_16_rsp_i_ack, dev_16_rsp_i_data};
  assign n1864_o = n1924_o[31:0]; // extract
  assign n1865_o = n1924_o[63:32]; // extract
  assign n1866_o = n1924_o[67:64]; // extract
  assign n1867_o = n1924_o[68]; // extract
  assign n1868_o = n1924_o[69]; // extract
  assign n1869_o = n1924_o[70]; // extract
  assign n1870_o = n1924_o[71]; // extract
  assign n1871_o = n1924_o[72]; // extract
  assign n1872_o = n1924_o[73]; // extract
  assign n1873_o = {dev_17_rsp_i_err, dev_17_rsp_i_ack, dev_17_rsp_i_data};
  assign n1875_o = n1925_o[31:0]; // extract
  assign n1876_o = n1925_o[63:32]; // extract
  assign n1877_o = n1925_o[67:64]; // extract
  assign n1878_o = n1925_o[68]; // extract
  assign n1879_o = n1925_o[69]; // extract
  assign n1880_o = n1925_o[70]; // extract
  assign n1881_o = n1925_o[71]; // extract
  assign n1882_o = n1925_o[72]; // extract
  assign n1883_o = n1925_o[73]; // extract
  assign n1884_o = {dev_18_rsp_i_err, dev_18_rsp_i_ack, dev_18_rsp_i_data};
  assign n1886_o = n1926_o[31:0]; // extract
  assign n1887_o = n1926_o[63:32]; // extract
  assign n1888_o = n1926_o[67:64]; // extract
  assign n1889_o = n1926_o[68]; // extract
  assign n1890_o = n1926_o[69]; // extract
  assign n1891_o = n1926_o[70]; // extract
  assign n1892_o = n1926_o[71]; // extract
  assign n1893_o = n1926_o[72]; // extract
  assign n1894_o = n1926_o[73]; // extract
  assign n1895_o = {dev_19_rsp_i_err, dev_19_rsp_i_ack, dev_19_rsp_i_data};
  assign n1897_o = n1927_o[31:0]; // extract
  assign n1898_o = n1927_o[63:32]; // extract
  assign n1899_o = n1927_o[67:64]; // extract
  assign n1900_o = n1927_o[68]; // extract
  assign n1901_o = n1927_o[69]; // extract
  assign n1902_o = n1927_o[70]; // extract
  assign n1903_o = n1927_o[71]; // extract
  assign n1904_o = n1927_o[72]; // extract
  assign n1905_o = n1927_o[73]; // extract
  assign n1906_o = {dev_20_rsp_i_err, dev_20_rsp_i_ack, dev_20_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:532:10  */
  assign dev_req = n1987_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:533:10  */
  assign dev_rsp = n1988_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:539:26  */
  assign n1907_o = dev_req[1553:1480]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:540:26  */
  assign n1908_o = dev_req[1479:1406]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:541:26  */
  assign n1909_o = dev_req[1405:1332]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:542:26  */
  assign n1910_o = dev_req[1331:1258]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:543:26  */
  assign n1911_o = dev_req[1257:1184]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:544:26  */
  assign n1912_o = dev_req[1183:1110]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:545:26  */
  assign n1913_o = dev_req[1109:1036]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:546:26  */
  assign n1914_o = dev_req[1035:962]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:547:26  */
  assign n1915_o = dev_req[961:888]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:548:26  */
  assign n1916_o = dev_req[887:814]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:549:26  */
  assign n1917_o = dev_req[813:740]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:550:26  */
  assign n1918_o = dev_req[739:666]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:551:26  */
  assign n1919_o = dev_req[665:592]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:552:26  */
  assign n1920_o = dev_req[591:518]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:553:26  */
  assign n1921_o = dev_req[517:444]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:554:26  */
  assign n1922_o = dev_req[443:370]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:555:26  */
  assign n1923_o = dev_req[369:296]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:556:26  */
  assign n1924_o = dev_req[295:222]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:557:26  */
  assign n1925_o = dev_req[221:148]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:558:26  */
  assign n1926_o = dev_req[147:74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:559:26  */
  assign n1927_o = dev_req[73:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:572:28  */
  assign n1930_o = n1671_o[12:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:572:55  */
  assign n1932_o = n1930_o == 5'b11110;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:573:40  */
  assign n1933_o = n1671_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:572:9  */
  assign n1935_o = n1932_o ? n1933_o : 1'b0;
  assign n1936_o = n1671_o[73:69]; // extract
  assign n1937_o = n1671_o[67:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:572:28  */
  assign n1940_o = n1671_o[12:8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:572:55  */
  assign n1942_o = n1940_o == 5'b10100;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:573:40  */
  assign n1943_o = n1671_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:572:9  */
  assign n1945_o = n1942_o ? n1943_o : 1'b0;
  assign n1946_o = n1671_o[73:69]; // extract
  assign n1947_o = n1671_o[67:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:596:29  */
  assign n1952_o = n1951_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:596:48  */
  assign n1954_o = dev_rsp[677:646]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:596:34  */
  assign n1955_o = n1952_o | n1954_o;
  assign n1957_o = n1956_o[33:32]; // extract
  assign n1958_o = {n1957_o, n1955_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:597:29  */
  assign n1959_o = n1958_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:597:48  */
  assign n1961_o = dev_rsp[678]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:597:34  */
  assign n1962_o = n1959_o | n1961_o;
  assign n1963_o = n1956_o[33]; // extract
  assign n1964_o = {n1963_o, n1962_o, n1955_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:598:29  */
  assign n1965_o = n1964_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:598:48  */
  assign n1967_o = dev_rsp[679]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:598:34  */
  assign n1968_o = n1965_o | n1967_o;
  assign n1969_o = {n1968_o, n1962_o, n1955_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:596:29  */
  assign n1970_o = n1969_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:596:48  */
  assign n1972_o = dev_rsp[337:306]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:596:34  */
  assign n1973_o = n1970_o | n1972_o;
  assign n1974_o = {n1968_o, n1962_o, n1973_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:597:29  */
  assign n1975_o = n1974_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:597:48  */
  assign n1977_o = dev_rsp[338]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:597:34  */
  assign n1978_o = n1975_o | n1977_o;
  assign n1979_o = {n1968_o, n1978_o, n1973_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:598:29  */
  assign n1980_o = n1979_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:598:48  */
  assign n1982_o = dev_rsp[339]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:598:34  */
  assign n1983_o = n1980_o | n1982_o;
  assign n1984_o = {n1983_o, n1978_o, n1973_o};
  assign n1987_o = {74'b00000000000000000000000000000000000000000000000000000000000000000000000000, n1936_o, n1935_o, n1937_o, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, n1946_o, n1945_o, n1947_o, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000};
  assign n1988_o = {n1686_o, n1697_o, n1708_o, n1719_o, n1730_o, n1741_o, n1752_o, n1763_o, n1774_o, n1785_o, n1796_o, n1807_o, n1818_o, n1829_o, n1840_o, n1851_o, n1862_o, n1873_o, n1884_o, n1895_o, n1906_o};
endmodule

module neorv32_cache_32_32_b2a9daee4605f0af85049a2738d2ab5c0686fc65
  (input  clk_i,
   input  rstn_i,
   input  [31:0] host_req_i_addr,
   input  [31:0] host_req_i_data,
   input  [3:0] host_req_i_ben,
   input  host_req_i_stb,
   input  host_req_i_rw,
   input  host_req_i_src,
   input  host_req_i_priv,
   input  host_req_i_rvso,
   input  host_req_i_fence,
   input  [31:0] bus_rsp_i_data,
   input  bus_rsp_i_ack,
   input  bus_rsp_i_err,
   output [31:0] host_rsp_o_data,
   output host_rsp_o_ack,
   output host_rsp_o_err,
   output [31:0] bus_req_o_addr,
   output [31:0] bus_req_o_data,
   output [3:0] bus_req_o_ben,
   output bus_req_o_stb,
   output bus_req_o_rw,
   output bus_req_o_src,
   output bus_req_o_priv,
   output bus_req_o_rvso,
   output bus_req_o_fence);
  wire [73:0] n1468_o;
  wire [31:0] n1470_o;
  wire n1471_o;
  wire n1472_o;
  wire [31:0] n1474_o;
  wire [31:0] n1475_o;
  wire [3:0] n1476_o;
  wire n1477_o;
  wire n1478_o;
  wire n1479_o;
  wire n1480_o;
  wire n1481_o;
  wire n1482_o;
  wire [33:0] n1483_o;
  wire dir_acc_d;
  wire dir_acc_q;
  wire [73:0] bus_req;
  wire [73:0] dir_req_d;
  wire [73:0] dir_req_q;
  wire [73:0] cache_req;
  wire [33:0] bus_rsp;
  wire [33:0] dir_rsp_d;
  wire [33:0] dir_rsp_q;
  wire [33:0] cache_rsp;
  wire [69:0] cache_in_host;
  wire [69:0] cache_in_bus;
  wire [69:0] cache_in;
  wire [32:0] cache_out;
  wire cache_stat_dirty;
  wire cache_stat_hit;
  wire [31:0] cache_stat_base;
  wire cache_cmd_inval;
  wire cache_cmd_new;
  wire cache_cmd_dirty;
  wire bus_cmd_sync;
  wire bus_cmd_miss;
  wire bus_cmd_busy;
  wire [3:0] n1485_o;
  wire n1487_o;
  wire n1488_o;
  wire n1489_o;
  wire n1491_o;
  wire n1492_o;
  wire n1495_o;
  wire n1496_o;
  wire [67:0] n1498_o;
  wire [3:0] n1500_o;
  wire n1501_o;
  wire n1502_o;
  wire n1503_o;
  wire [4:0] n1504_o;
  wire [67:0] n1505_o;
  wire n1508_o;
  wire n1510_o;
  wire n1511_o;
  wire n1512_o;
  wire n1513_o;
  wire n1514_o;
  wire n1515_o;
  wire n1516_o;
  wire n1517_o;
  wire n1519_o;
  wire n1521_o;
  wire n1532_o;
  wire [33:0] n1533_o;
  wire [33:0] neorv32_cache_host_inst_n1534;
  wire neorv32_cache_host_inst_n1535;
  wire neorv32_cache_host_inst_n1536;
  wire neorv32_cache_host_inst_n1537;
  wire [31:0] neorv32_cache_host_inst_n1538;
  wire [3:0] neorv32_cache_host_inst_n1539;
  wire neorv32_cache_host_inst_n1540;
  wire [31:0] neorv32_cache_host_inst_n1541;
  wire neorv32_cache_host_inst_n1542;
  wire [31:0] n1543_o;
  wire n1544_o;
  wire [31:0] neorv32_cache_host_inst_rsp_o_data;
  wire neorv32_cache_host_inst_rsp_o_ack;
  wire neorv32_cache_host_inst_rsp_o_err;
  wire neorv32_cache_host_inst_bus_sync_o;
  wire neorv32_cache_host_inst_bus_miss_o;
  wire neorv32_cache_host_inst_dirty_o;
  wire [31:0] neorv32_cache_host_inst_addr_o;
  wire [3:0] neorv32_cache_host_inst_we_o;
  wire neorv32_cache_host_inst_swe_o;
  wire [31:0] neorv32_cache_host_inst_wdata_o;
  wire neorv32_cache_host_inst_wstat_o;
  wire [31:0] n1545_o;
  wire [31:0] n1546_o;
  wire [3:0] n1547_o;
  wire n1548_o;
  wire n1549_o;
  wire n1550_o;
  wire n1551_o;
  wire n1552_o;
  wire n1553_o;
  wire [33:0] n1554_o;
  wire neorv32_cache_memory_inst_n1573;
  wire neorv32_cache_memory_inst_n1574;
  wire [31:0] neorv32_cache_memory_inst_n1575;
  wire [31:0] n1576_o;
  wire [3:0] n1577_o;
  wire n1578_o;
  wire [31:0] n1579_o;
  wire n1580_o;
  wire [31:0] neorv32_cache_memory_inst_n1581;
  wire neorv32_cache_memory_inst_n1582;
  wire neorv32_cache_memory_inst_hit_o;
  wire neorv32_cache_memory_inst_dirty_o;
  wire [31:0] neorv32_cache_memory_inst_base_o;
  wire [31:0] neorv32_cache_memory_inst_rdata_o;
  wire neorv32_cache_memory_inst_rstat_o;
  wire n1593_o;
  wire [69:0] n1594_o;
  wire [73:0] neorv32_cache_bus_inst_n1595;
  wire neorv32_cache_bus_inst_n1596;
  wire neorv32_cache_bus_inst_n1597;
  wire neorv32_cache_bus_inst_n1598;
  wire [31:0] neorv32_cache_bus_inst_n1599;
  wire [3:0] neorv32_cache_bus_inst_n1600;
  wire neorv32_cache_bus_inst_n1601;
  wire [31:0] neorv32_cache_bus_inst_n1602;
  wire neorv32_cache_bus_inst_n1603;
  wire [31:0] n1604_o;
  wire [31:0] neorv32_cache_bus_inst_bus_req_o_addr;
  wire [31:0] neorv32_cache_bus_inst_bus_req_o_data;
  wire [3:0] neorv32_cache_bus_inst_bus_req_o_ben;
  wire neorv32_cache_bus_inst_bus_req_o_stb;
  wire neorv32_cache_bus_inst_bus_req_o_rw;
  wire neorv32_cache_bus_inst_bus_req_o_src;
  wire neorv32_cache_bus_inst_bus_req_o_priv;
  wire neorv32_cache_bus_inst_bus_req_o_rvso;
  wire neorv32_cache_bus_inst_bus_req_o_fence;
  wire neorv32_cache_bus_inst_cmd_busy_o;
  wire neorv32_cache_bus_inst_inval_o;
  wire neorv32_cache_bus_inst_new_o;
  wire [31:0] neorv32_cache_bus_inst_addr_o;
  wire [3:0] neorv32_cache_bus_inst_we_o;
  wire neorv32_cache_bus_inst_swe_o;
  wire [31:0] neorv32_cache_bus_inst_wdata_o;
  wire neorv32_cache_bus_inst_wstat_o;
  wire [31:0] n1605_o;
  wire [31:0] n1606_o;
  wire [3:0] n1607_o;
  wire n1608_o;
  wire n1609_o;
  wire n1610_o;
  wire n1611_o;
  wire n1612_o;
  wire n1613_o;
  wire [73:0] n1614_o;
  wire [31:0] n1616_o;
  wire n1617_o;
  wire n1618_o;
  wire [31:0] bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_data;
  wire bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_ack;
  wire bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_err;
  wire [31:0] bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_data;
  wire bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_ack;
  wire bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_err;
  wire [31:0] bus_switch_enable_neorv32_cache_bus_switch_x_req_o_addr;
  wire [31:0] bus_switch_enable_neorv32_cache_bus_switch_x_req_o_data;
  wire [3:0] bus_switch_enable_neorv32_cache_bus_switch_x_req_o_ben;
  wire bus_switch_enable_neorv32_cache_bus_switch_x_req_o_stb;
  wire bus_switch_enable_neorv32_cache_bus_switch_x_req_o_rw;
  wire bus_switch_enable_neorv32_cache_bus_switch_x_req_o_src;
  wire bus_switch_enable_neorv32_cache_bus_switch_x_req_o_priv;
  wire bus_switch_enable_neorv32_cache_bus_switch_x_req_o_rvso;
  wire bus_switch_enable_neorv32_cache_bus_switch_x_req_o_fence;
  wire [31:0] n1636_o;
  wire [31:0] n1637_o;
  wire [3:0] n1638_o;
  wire n1639_o;
  wire n1640_o;
  wire n1641_o;
  wire n1642_o;
  wire n1643_o;
  wire n1644_o;
  wire [33:0] n1645_o;
  wire [31:0] n1647_o;
  wire [31:0] n1648_o;
  wire [3:0] n1649_o;
  wire n1650_o;
  wire n1651_o;
  wire n1652_o;
  wire n1653_o;
  wire n1654_o;
  wire n1655_o;
  wire [33:0] n1656_o;
  wire [73:0] n1658_o;
  wire [31:0] n1660_o;
  wire n1661_o;
  wire n1662_o;
  reg n1663_q;
  wire [73:0] n1664_o;
  reg [73:0] n1665_q;
  wire [73:0] n1666_o;
  reg [33:0] n1667_q;
  wire [69:0] n1668_o;
  wire [69:0] n1669_o;
  wire [32:0] n1670_o;
  assign host_rsp_o_data = n1470_o; //(module output)
  assign host_rsp_o_ack = n1471_o; //(module output)
  assign host_rsp_o_err = n1472_o; //(module output)
  assign bus_req_o_addr = n1474_o; //(module output)
  assign bus_req_o_data = n1475_o; //(module output)
  assign bus_req_o_ben = n1476_o; //(module output)
  assign bus_req_o_stb = n1477_o; //(module output)
  assign bus_req_o_rw = n1478_o; //(module output)
  assign bus_req_o_src = n1479_o; //(module output)
  assign bus_req_o_priv = n1480_o; //(module output)
  assign bus_req_o_rvso = n1481_o; //(module output)
  assign bus_req_o_fence = n1482_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:67:5  */
  assign n1468_o = {host_req_i_fence, host_req_i_rvso, host_req_i_priv, host_req_i_src, host_req_i_rw, host_req_i_stb, host_req_i_ben, host_req_i_data, host_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:65:5  */
  assign n1470_o = n1533_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:64:5  */
  assign n1471_o = n1533_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:62:5  */
  assign n1472_o = n1533_o[33]; // extract
  assign n1474_o = n1658_o[31:0]; // extract
  assign n1475_o = n1658_o[63:32]; // extract
  assign n1476_o = n1658_o[67:64]; // extract
  assign n1477_o = n1658_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1022:14  */
  assign n1478_o = n1658_o[69]; // extract
  assign n1479_o = n1658_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:716:12  */
  assign n1480_o = n1658_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:716:12  */
  assign n1481_o = n1658_o[72]; // extract
  assign n1482_o = n1658_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:716:12  */
  assign n1483_o = {bus_rsp_i_err, bus_rsp_i_ack, bus_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:172:10  */
  assign dir_acc_d = n1492_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:172:21  */
  assign dir_acc_q = n1663_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:175:10  */
  assign bus_req = neorv32_cache_bus_inst_n1595; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:175:19  */
  assign dir_req_d = n1664_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:175:30  */
  assign dir_req_q = n1665_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:175:41  */
  assign cache_req = n1666_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:176:10  */
  assign bus_rsp = n1645_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:176:19  */
  assign dir_rsp_d = n1656_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:176:30  */
  assign dir_rsp_q = n1667_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:176:41  */
  assign cache_rsp = neorv32_cache_host_inst_n1534; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:186:10  */
  assign cache_in_host = n1668_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:186:25  */
  assign cache_in_bus = n1669_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:186:39  */
  assign cache_in = n1594_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:192:10  */
  assign cache_out = n1670_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:195:10  */
  assign cache_stat_dirty = neorv32_cache_memory_inst_n1574; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:195:28  */
  assign cache_stat_hit = neorv32_cache_memory_inst_n1573; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:196:10  */
  assign cache_stat_base = neorv32_cache_memory_inst_n1575; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:199:10  */
  assign cache_cmd_inval = neorv32_cache_bus_inst_n1597; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:199:27  */
  assign cache_cmd_new = neorv32_cache_bus_inst_n1598; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:199:42  */
  assign cache_cmd_dirty = neorv32_cache_host_inst_n1537; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:199:59  */
  assign bus_cmd_sync = neorv32_cache_host_inst_n1535; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:199:73  */
  assign bus_cmd_miss = neorv32_cache_host_inst_n1536; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:199:87  */
  assign bus_cmd_busy = neorv32_cache_bus_inst_n1596; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:206:42  */
  assign n1485_o = n1468_o[31:28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:206:57  */
  assign n1487_o = $unsigned(n1485_o) >= $unsigned(4'b1111);
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:207:38  */
  assign n1488_o = n1468_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:206:70  */
  assign n1489_o = n1487_o | n1488_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:205:44  */
  assign n1491_o = n1489_o & 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:205:20  */
  assign n1492_o = n1491_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:216:35  */
  assign n1495_o = n1468_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:216:39  */
  assign n1496_o = n1495_o & dir_acc_d;
  assign n1498_o = n1468_o[67:0]; // extract
  assign n1500_o = n1468_o[72:69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:219:33  */
  assign n1501_o = n1468_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:219:42  */
  assign n1502_o = ~dir_acc_d;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:219:37  */
  assign n1503_o = n1501_o & n1502_o;
  assign n1504_o = n1468_o[73:69]; // extract
  assign n1505_o = n1468_o[67:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:227:18  */
  assign n1508_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:232:23  */
  assign n1510_o = ~dir_acc_q;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:232:46  */
  assign n1511_o = n1468_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:232:30  */
  assign n1512_o = n1511_o & n1510_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:232:57  */
  assign n1513_o = dir_acc_d & n1512_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:234:49  */
  assign n1514_o = dir_rsp_q[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:234:74  */
  assign n1515_o = dir_rsp_q[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:234:60  */
  assign n1516_o = n1514_o | n1515_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:234:33  */
  assign n1517_o = n1516_o & dir_acc_q;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:234:9  */
  assign n1519_o = n1517_o ? 1'b0 : dir_acc_q;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:232:9  */
  assign n1521_o = n1513_o ? 1'b1 : n1519_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:250:45  */
  assign n1532_o = ~dir_acc_q;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:250:29  */
  assign n1533_o = n1532_o ? cache_rsp : dir_rsp_q;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:275:19  */
  assign neorv32_cache_host_inst_n1534 = n1554_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:277:19  */
  assign neorv32_cache_host_inst_n1535 = neorv32_cache_host_inst_bus_sync_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:278:19  */
  assign neorv32_cache_host_inst_n1536 = neorv32_cache_host_inst_bus_miss_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:281:19  */
  assign neorv32_cache_host_inst_n1537 = neorv32_cache_host_inst_dirty_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:284:19  */
  assign neorv32_cache_host_inst_n1538 = neorv32_cache_host_inst_addr_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:285:19  */
  assign neorv32_cache_host_inst_n1539 = neorv32_cache_host_inst_we_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:286:19  */
  assign neorv32_cache_host_inst_n1540 = neorv32_cache_host_inst_swe_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:287:19  */
  assign neorv32_cache_host_inst_n1541 = neorv32_cache_host_inst_wdata_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:288:19  */
  assign neorv32_cache_host_inst_n1542 = neorv32_cache_host_inst_wstat_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:289:29  */
  assign n1543_o = cache_out[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:290:29  */
  assign n1544_o = cache_out[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:265:3  */
  neorv32_cache_host_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_cache_host_inst (
    .rstn_i(rstn_i),
    .clk_i(clk_i),
    .req_i_addr(n1545_o),
    .req_i_data(n1546_o),
    .req_i_ben(n1547_o),
    .req_i_stb(n1548_o),
    .req_i_rw(n1549_o),
    .req_i_src(n1550_o),
    .req_i_priv(n1551_o),
    .req_i_rvso(n1552_o),
    .req_i_fence(n1553_o),
    .bus_busy_i(bus_cmd_busy),
    .hit_i(cache_stat_hit),
    .rdata_i(n1543_o),
    .rstat_i(n1544_o),
    .rsp_o_data(neorv32_cache_host_inst_rsp_o_data),
    .rsp_o_ack(neorv32_cache_host_inst_rsp_o_ack),
    .rsp_o_err(neorv32_cache_host_inst_rsp_o_err),
    .bus_sync_o(neorv32_cache_host_inst_bus_sync_o),
    .bus_miss_o(neorv32_cache_host_inst_bus_miss_o),
    .dirty_o(neorv32_cache_host_inst_dirty_o),
    .addr_o(neorv32_cache_host_inst_addr_o),
    .we_o(neorv32_cache_host_inst_we_o),
    .swe_o(neorv32_cache_host_inst_swe_o),
    .wdata_o(neorv32_cache_host_inst_wdata_o),
    .wstat_o(neorv32_cache_host_inst_wstat_o));
  assign n1545_o = cache_req[31:0]; // extract
  assign n1546_o = cache_req[63:32]; // extract
  assign n1547_o = cache_req[67:64]; // extract
  assign n1548_o = cache_req[68]; // extract
  assign n1549_o = cache_req[69]; // extract
  assign n1550_o = cache_req[70]; // extract
  assign n1551_o = cache_req[71]; // extract
  assign n1552_o = cache_req[72]; // extract
  assign n1553_o = cache_req[73]; // extract
  assign n1554_o = {neorv32_cache_host_inst_rsp_o_err, neorv32_cache_host_inst_rsp_o_ack, neorv32_cache_host_inst_rsp_o_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:311:17  */
  assign neorv32_cache_memory_inst_n1573 = neorv32_cache_memory_inst_hit_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:312:17  */
  assign neorv32_cache_memory_inst_n1574 = neorv32_cache_memory_inst_dirty_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:313:17  */
  assign neorv32_cache_memory_inst_n1575 = neorv32_cache_memory_inst_base_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:315:26  */
  assign n1576_o = cache_in[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:316:26  */
  assign n1577_o = cache_in[35:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:317:26  */
  assign n1578_o = cache_in[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:318:26  */
  assign n1579_o = cache_in[68:37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:319:26  */
  assign n1580_o = cache_in[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:320:17  */
  assign neorv32_cache_memory_inst_n1581 = neorv32_cache_memory_inst_rdata_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:321:17  */
  assign neorv32_cache_memory_inst_n1582 = neorv32_cache_memory_inst_rstat_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:296:3  */
  neorv32_cache_memory_32_32_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_cache_memory_inst (
    .rstn_i(rstn_i),
    .clk_i(clk_i),
    .inval_i(cache_cmd_inval),
    .new_i(cache_cmd_new),
    .dirty_i(cache_cmd_dirty),
    .addr_i(n1576_o),
    .we_i(n1577_o),
    .swe_i(n1578_o),
    .wdata_i(n1579_o),
    .wstat_i(n1580_o),
    .hit_o(neorv32_cache_memory_inst_hit_o),
    .dirty_o(neorv32_cache_memory_inst_dirty_o),
    .base_o(neorv32_cache_memory_inst_base_o),
    .rdata_o(neorv32_cache_memory_inst_rdata_o),
    .rstat_o(neorv32_cache_memory_inst_rstat_o));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:325:48  */
  assign n1593_o = ~bus_cmd_busy;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:325:29  */
  assign n1594_o = n1593_o ? cache_in_host : cache_in_bus;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:343:19  */
  assign neorv32_cache_bus_inst_n1595 = n1614_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:348:19  */
  assign neorv32_cache_bus_inst_n1596 = neorv32_cache_bus_inst_cmd_busy_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:350:19  */
  assign neorv32_cache_bus_inst_n1597 = neorv32_cache_bus_inst_inval_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:351:19  */
  assign neorv32_cache_bus_inst_n1598 = neorv32_cache_bus_inst_new_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:355:19  */
  assign neorv32_cache_bus_inst_n1599 = neorv32_cache_bus_inst_addr_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:356:19  */
  assign neorv32_cache_bus_inst_n1600 = neorv32_cache_bus_inst_we_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:357:19  */
  assign neorv32_cache_bus_inst_n1601 = neorv32_cache_bus_inst_swe_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:358:19  */
  assign neorv32_cache_bus_inst_n1602 = neorv32_cache_bus_inst_wdata_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:359:19  */
  assign neorv32_cache_bus_inst_n1603 = neorv32_cache_bus_inst_wstat_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:360:29  */
  assign n1604_o = cache_out[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:330:3  */
  neorv32_cache_bus_32_32_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_cache_bus_inst (
    .rstn_i(rstn_i),
    .clk_i(clk_i),
    .host_req_i_addr(n1605_o),
    .host_req_i_data(n1606_o),
    .host_req_i_ben(n1607_o),
    .host_req_i_stb(n1608_o),
    .host_req_i_rw(n1609_o),
    .host_req_i_src(n1610_o),
    .host_req_i_priv(n1611_o),
    .host_req_i_rvso(n1612_o),
    .host_req_i_fence(n1613_o),
    .bus_rsp_i_data(n1616_o),
    .bus_rsp_i_ack(n1617_o),
    .bus_rsp_i_err(n1618_o),
    .cmd_sync_i(bus_cmd_sync),
    .cmd_miss_i(bus_cmd_miss),
    .dirty_i(cache_stat_dirty),
    .base_i(cache_stat_base),
    .rdata_i(n1604_o),
    .bus_req_o_addr(neorv32_cache_bus_inst_bus_req_o_addr),
    .bus_req_o_data(neorv32_cache_bus_inst_bus_req_o_data),
    .bus_req_o_ben(neorv32_cache_bus_inst_bus_req_o_ben),
    .bus_req_o_stb(neorv32_cache_bus_inst_bus_req_o_stb),
    .bus_req_o_rw(neorv32_cache_bus_inst_bus_req_o_rw),
    .bus_req_o_src(neorv32_cache_bus_inst_bus_req_o_src),
    .bus_req_o_priv(neorv32_cache_bus_inst_bus_req_o_priv),
    .bus_req_o_rvso(neorv32_cache_bus_inst_bus_req_o_rvso),
    .bus_req_o_fence(neorv32_cache_bus_inst_bus_req_o_fence),
    .cmd_busy_o(neorv32_cache_bus_inst_cmd_busy_o),
    .inval_o(neorv32_cache_bus_inst_inval_o),
    .new_o(neorv32_cache_bus_inst_new_o),
    .addr_o(neorv32_cache_bus_inst_addr_o),
    .we_o(neorv32_cache_bus_inst_we_o),
    .swe_o(neorv32_cache_bus_inst_swe_o),
    .wdata_o(neorv32_cache_bus_inst_wdata_o),
    .wstat_o(neorv32_cache_bus_inst_wstat_o));
  assign n1605_o = n1468_o[31:0]; // extract
  assign n1606_o = n1468_o[63:32]; // extract
  assign n1607_o = n1468_o[67:64]; // extract
  assign n1608_o = n1468_o[68]; // extract
  assign n1609_o = n1468_o[69]; // extract
  assign n1610_o = n1468_o[70]; // extract
  assign n1611_o = n1468_o[71]; // extract
  assign n1612_o = n1468_o[72]; // extract
  assign n1613_o = n1468_o[73]; // extract
  assign n1614_o = {neorv32_cache_bus_inst_bus_req_o_fence, neorv32_cache_bus_inst_bus_req_o_rvso, neorv32_cache_bus_inst_bus_req_o_priv, neorv32_cache_bus_inst_bus_req_o_src, neorv32_cache_bus_inst_bus_req_o_rw, neorv32_cache_bus_inst_bus_req_o_stb, neorv32_cache_bus_inst_bus_req_o_ben, neorv32_cache_bus_inst_bus_req_o_data, neorv32_cache_bus_inst_bus_req_o_addr};
  assign n1616_o = bus_rsp[31:0]; // extract
  assign n1617_o = bus_rsp[32]; // extract
  assign n1618_o = bus_rsp[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:370:5  */
  neorv32_bus_switch_1489f923c4dca729178b3e3233458550d8dddf29 bus_switch_enable_neorv32_cache_bus_switch (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .a_req_i_addr(n1636_o),
    .a_req_i_data(n1637_o),
    .a_req_i_ben(n1638_o),
    .a_req_i_stb(n1639_o),
    .a_req_i_rw(n1640_o),
    .a_req_i_src(n1641_o),
    .a_req_i_priv(n1642_o),
    .a_req_i_rvso(n1643_o),
    .a_req_i_fence(n1644_o),
    .b_req_i_addr(n1647_o),
    .b_req_i_data(n1648_o),
    .b_req_i_ben(n1649_o),
    .b_req_i_stb(n1650_o),
    .b_req_i_rw(n1651_o),
    .b_req_i_src(n1652_o),
    .b_req_i_priv(n1653_o),
    .b_req_i_rvso(n1654_o),
    .b_req_i_fence(n1655_o),
    .x_rsp_i_data(n1660_o),
    .x_rsp_i_ack(n1661_o),
    .x_rsp_i_err(n1662_o),
    .a_rsp_o_data(bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_data),
    .a_rsp_o_ack(bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_ack),
    .a_rsp_o_err(bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_err),
    .b_rsp_o_data(bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_data),
    .b_rsp_o_ack(bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_ack),
    .b_rsp_o_err(bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_err),
    .x_req_o_addr(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_addr),
    .x_req_o_data(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_data),
    .x_req_o_ben(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_ben),
    .x_req_o_stb(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_stb),
    .x_req_o_rw(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_rw),
    .x_req_o_src(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_src),
    .x_req_o_priv(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_priv),
    .x_req_o_rvso(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_rvso),
    .x_req_o_fence(bus_switch_enable_neorv32_cache_bus_switch_x_req_o_fence));
  assign n1636_o = bus_req[31:0]; // extract
  assign n1637_o = bus_req[63:32]; // extract
  assign n1638_o = bus_req[67:64]; // extract
  assign n1639_o = bus_req[68]; // extract
  assign n1640_o = bus_req[69]; // extract
  assign n1641_o = bus_req[70]; // extract
  assign n1642_o = bus_req[71]; // extract
  assign n1643_o = bus_req[72]; // extract
  assign n1644_o = bus_req[73]; // extract
  assign n1645_o = {bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_err, bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_ack, bus_switch_enable_neorv32_cache_bus_switch_a_rsp_o_data};
  assign n1647_o = dir_req_q[31:0]; // extract
  assign n1648_o = dir_req_q[63:32]; // extract
  assign n1649_o = dir_req_q[67:64]; // extract
  assign n1650_o = dir_req_q[68]; // extract
  assign n1651_o = dir_req_q[69]; // extract
  assign n1652_o = dir_req_q[70]; // extract
  assign n1653_o = dir_req_q[71]; // extract
  assign n1654_o = dir_req_q[72]; // extract
  assign n1655_o = dir_req_q[73]; // extract
  assign n1656_o = {bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_err, bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_ack, bus_switch_enable_neorv32_cache_bus_switch_b_rsp_o_data};
  assign n1658_o = {bus_switch_enable_neorv32_cache_bus_switch_x_req_o_fence, bus_switch_enable_neorv32_cache_bus_switch_x_req_o_rvso, bus_switch_enable_neorv32_cache_bus_switch_x_req_o_priv, bus_switch_enable_neorv32_cache_bus_switch_x_req_o_src, bus_switch_enable_neorv32_cache_bus_switch_x_req_o_rw, bus_switch_enable_neorv32_cache_bus_switch_x_req_o_stb, bus_switch_enable_neorv32_cache_bus_switch_x_req_o_ben, bus_switch_enable_neorv32_cache_bus_switch_x_req_o_data, bus_switch_enable_neorv32_cache_bus_switch_x_req_o_addr};
  assign n1660_o = n1483_o[31:0]; // extract
  assign n1661_o = n1483_o[32]; // extract
  assign n1662_o = n1483_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:231:7  */
  always @(posedge clk_i or posedge n1508_o)
    if (n1508_o)
      n1663_q <= 1'b0;
    else
      n1663_q <= n1521_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:227:7  */
  assign n1664_o = {1'b0, n1500_o, n1496_o, n1498_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:231:7  */
  always @(posedge clk_i or posedge n1508_o)
    if (n1508_o)
      n1665_q <= 74'b00000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n1665_q <= dir_req_d;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:227:7  */
  assign n1666_o = {n1504_o, n1503_o, n1505_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:231:7  */
  always @(posedge clk_i or posedge n1508_o)
    if (n1508_o)
      n1667_q <= 34'b0000000000000000000000000000000000;
    else
      n1667_q <= dir_rsp_d;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cache.vhd:227:7  */
  assign n1668_o = {neorv32_cache_host_inst_n1542, neorv32_cache_host_inst_n1541, neorv32_cache_host_inst_n1540, neorv32_cache_host_inst_n1539, neorv32_cache_host_inst_n1538};
  assign n1669_o = {neorv32_cache_bus_inst_n1603, neorv32_cache_bus_inst_n1602, neorv32_cache_bus_inst_n1601, neorv32_cache_bus_inst_n1600, neorv32_cache_bus_inst_n1599};
  assign n1670_o = {neorv32_cache_memory_inst_n1582, neorv32_cache_memory_inst_n1581};
endmodule

module neorv32_xbus_1024_eee447edc79fea1ca7c7d34e463261cda4ba339e
  (input  clk_i,
   input  rstn_i,
   input  [31:0] bus_req_i_addr,
   input  [31:0] bus_req_i_data,
   input  [3:0] bus_req_i_ben,
   input  bus_req_i_stb,
   input  bus_req_i_rw,
   input  bus_req_i_src,
   input  bus_req_i_priv,
   input  bus_req_i_rvso,
   input  bus_req_i_fence,
   input  [31:0] xbus_dat_i,
   input  xbus_ack_i,
   input  xbus_err_i,
   output [31:0] bus_rsp_o_data,
   output bus_rsp_o_ack,
   output bus_rsp_o_err,
   output [31:0] xbus_adr_o,
   output [31:0] xbus_dat_o,
   output xbus_we_o,
   output [3:0] xbus_sel_o,
   output xbus_stb_o,
   output xbus_cyc_o);
  wire [73:0] n1300_o;
  wire [31:0] n1302_o;
  wire n1303_o;
  wire n1304_o;
  wire [115:0] ctrl;
  wire stb_int;
  wire cyc_int;
  wire ack_gated;
  wire err_gated;
  wire [31:0] rdata_gated;
  wire n1316_o;
  wire n1328_o;
  wire n1334_o;
  wire n1335_o;
  wire n1336_o;
  wire n1337_o;
  wire [31:0] n1338_o;
  wire [31:0] n1339_o;
  wire [3:0] n1340_o;
  wire [64:0] n1342_o;
  wire n1343_o;
  wire n1344_o;
  wire [64:0] n1345_o;
  wire [64:0] n1346_o;
  wire [3:0] n1347_o;
  wire [3:0] n1348_o;
  wire n1349_o;
  wire n1350_o;
  wire [31:0] n1351_o;
  wire n1361_o;
  wire n1363_o;
  wire n1365_o;
  wire n1366_o;
  wire n1367_o;
  wire n1368_o;
  wire n1369_o;
  wire n1370_o;
  wire n1371_o;
  wire n1372_o;
  wire n1373_o;
  wire n1374_o;
  wire n1375_o;
  wire n1376_o;
  wire n1377_o;
  wire n1378_o;
  wire n1379_o;
  wire n1380_o;
  wire n1381_o;
  wire n1382_o;
  wire n1383_o;
  wire n1384_o;
  wire n1385_o;
  wire n1387_o;
  wire n1388_o;
  wire n1391_o;
  wire n1392_o;
  wire n1393_o;
  wire n1394_o;
  wire n1395_o;
  wire n1396_o;
  wire [10:0] n1397_o;
  wire [10:0] n1399_o;
  wire [12:0] n1400_o;
  wire n1401_o;
  wire n1403_o;
  wire [31:0] n1404_o;
  wire n1406_o;
  wire [12:0] n1407_o;
  wire [12:0] n1408_o;
  wire [115:0] n1409_o;
  wire [115:0] n1411_o;
  wire n1414_o;
  wire n1416_o;
  wire n1417_o;
  wire n1418_o;
  wire n1419_o;
  wire n1420_o;
  wire n1421_o;
  wire n1422_o;
  wire n1423_o;
  wire n1425_o;
  wire n1426_o;
  wire [31:0] n1427_o;
  wire [31:0] n1429_o;
  wire [31:0] n1430_o;
  wire [31:0] n1431_o;
  wire [31:0] n1433_o;
  wire [31:0] n1434_o;
  wire n1435_o;
  wire n1437_o;
  wire n1438_o;
  wire [3:0] n1439_o;
  wire [3:0] n1441_o;
  wire [3:0] n1442_o;
  wire n1444_o;
  wire n1445_o;
  wire n1446_o;
  wire n1448_o;
  wire n1449_o;
  wire n1451_o;
  wire n1452_o;
  wire n1453_o;
  wire n1454_o;
  wire [31:0] n1455_o;
  wire [31:0] n1457_o;
  wire [31:0] n1459_o;
  wire n1460_o;
  wire n1462_o;
  wire n1463_o;
  wire n1465_o;
  reg [115:0] n1466_q;
  wire [33:0] n1467_o;
  assign bus_rsp_o_data = n1302_o; //(module output)
  assign bus_rsp_o_ack = n1303_o; //(module output)
  assign bus_rsp_o_err = n1304_o; //(module output)
  assign xbus_adr_o = n1429_o; //(module output)
  assign xbus_dat_o = n1433_o; //(module output)
  assign xbus_we_o = n1437_o; //(module output)
  assign xbus_sel_o = n1441_o; //(module output)
  assign xbus_stb_o = n1444_o; //(module output)
  assign xbus_cyc_o = cyc_int; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:264:5  */
  assign n1300_o = {bus_req_i_fence, bus_req_i_rvso, bus_req_i_priv, bus_req_i_src, bus_req_i_rw, bus_req_i_stb, bus_req_i_ben, bus_req_i_data, bus_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:260:5  */
  assign n1302_o = n1467_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:258:5  */
  assign n1303_o = n1467_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:256:5  */
  assign n1304_o = n1467_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:95:10  */
  assign ctrl = n1466_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:96:10  */
  assign stb_int = n1416_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:97:10  */
  assign cyc_int = n1425_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:100:10  */
  assign ack_gated = n1446_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:101:10  */
  assign err_gated = n1449_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:102:10  */
  assign rdata_gated = n1455_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:129:16  */
  assign n1316_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:142:29  */
  assign n1328_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:16  */
  assign n1334_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:22  */
  assign n1335_o = ~n1334_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:150:23  */
  assign n1336_o = n1300_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:152:35  */
  assign n1337_o = n1300_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:153:35  */
  assign n1338_o = n1300_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:154:35  */
  assign n1339_o = n1300_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:155:35  */
  assign n1340_o = n1300_o[67:64]; // extract
  assign n1342_o = {n1339_o, n1338_o, n1337_o};
  assign n1343_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:150:9  */
  assign n1344_o = n1336_o ? 1'b1 : n1343_o;
  assign n1345_o = ctrl[66:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:7  */
  assign n1346_o = n1403_o ? n1342_o : n1345_o;
  assign n1347_o = ctrl[102:99]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:7  */
  assign n1348_o = n1406_o ? n1340_o : n1347_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:160:18  */
  assign n1349_o = ctrl[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:160:21  */
  assign n1350_o = ~n1349_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:160:9  */
  assign n1351_o = n1350_o ? xbus_dat_i : 32'b00000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1361_o = ctrl[115]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1363_o = 1'b0 | n1361_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1365_o = ctrl[114]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1366_o = n1363_o | n1365_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1367_o = ctrl[113]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1368_o = n1366_o | n1367_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1369_o = ctrl[112]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1370_o = n1368_o | n1369_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1371_o = ctrl[111]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1372_o = n1370_o | n1371_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1373_o = ctrl[110]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1374_o = n1372_o | n1373_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1375_o = ctrl[109]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1376_o = n1374_o | n1375_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1377_o = ctrl[108]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1378_o = n1376_o | n1377_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1379_o = ctrl[107]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1380_o = n1378_o | n1379_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1381_o = ctrl[106]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1382_o = n1380_o | n1381_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1383_o = ctrl[105]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1384_o = n1382_o | n1383_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:166:91  */
  assign n1385_o = ~n1384_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:166:60  */
  assign n1387_o = n1385_o & 1'b1;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:166:34  */
  assign n1388_o = xbus_err_i | n1387_o;
  assign n1391_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:166:9  */
  assign n1392_o = n1388_o ? 1'b0 : n1391_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:166:9  */
  assign n1393_o = n1388_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:163:9  */
  assign n1394_o = xbus_ack_i ? 1'b0 : n1392_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:163:9  */
  assign n1395_o = xbus_ack_i ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:163:9  */
  assign n1396_o = xbus_ack_i ? 1'b0 : n1393_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:172:59  */
  assign n1397_o = ctrl[115:105]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:172:68  */
  assign n1399_o = n1397_o - 11'b00000000001;
  assign n1400_o = {n1399_o, n1396_o, n1395_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:7  */
  assign n1401_o = n1335_o ? n1344_o : n1394_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:7  */
  assign n1403_o = n1336_o & n1335_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:7  */
  assign n1404_o = n1335_o ? 32'b00000000000000000000000000000000 : n1351_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:7  */
  assign n1406_o = n1336_o & n1335_o;
  assign n1407_o = {11'b10000000000, 1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:148:7  */
  assign n1408_o = n1335_o ? n1407_o : n1400_o;
  assign n1409_o = {n1408_o, n1348_o, n1404_o, n1346_o, n1328_o, n1401_o};
  assign n1411_o = {11'b00000000000, 1'b0, 1'b0, 4'b0000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 1'b0, 1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:179:25  */
  assign n1414_o = n1300_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:179:44  */
  assign n1416_o = 1'b1 ? n1414_o : n1420_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:179:78  */
  assign n1417_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:179:98  */
  assign n1418_o = ctrl[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:179:89  */
  assign n1419_o = ~n1418_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:179:84  */
  assign n1420_o = n1417_o & n1419_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:180:25  */
  assign n1421_o = n1300_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:180:37  */
  assign n1422_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:180:29  */
  assign n1423_o = n1421_o | n1422_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:180:44  */
  assign n1425_o = 1'b1 ? n1423_o : n1426_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:180:78  */
  assign n1426_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:182:27  */
  assign n1427_o = n1300_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:182:32  */
  assign n1429_o = 1'b1 ? n1427_o : n1430_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:182:66  */
  assign n1430_o = ctrl[34:3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:183:27  */
  assign n1431_o = n1300_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:183:32  */
  assign n1433_o = 1'b1 ? n1431_o : n1434_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:183:66  */
  assign n1434_o = ctrl[66:35]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:184:27  */
  assign n1435_o = n1300_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:184:32  */
  assign n1437_o = 1'b1 ? n1435_o : n1438_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:184:66  */
  assign n1438_o = ctrl[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:185:27  */
  assign n1439_o = n1300_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:185:32  */
  assign n1441_o = 1'b1 ? n1439_o : n1442_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:185:66  */
  assign n1442_o = ctrl[102:99]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:186:32  */
  assign n1444_o = 1'b0 ? stb_int : cyc_int;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:190:40  */
  assign n1445_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:190:29  */
  assign n1446_o = n1445_o ? xbus_ack_i : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:191:40  */
  assign n1448_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:191:29  */
  assign n1449_o = n1448_o ? xbus_err_i : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:192:40  */
  assign n1451_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:192:63  */
  assign n1452_o = ctrl[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:192:66  */
  assign n1453_o = ~n1452_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:192:53  */
  assign n1454_o = n1453_o & n1451_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:192:29  */
  assign n1455_o = n1454_o ? xbus_dat_i : 32'b00000000000000000000000000000000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:194:26  */
  assign n1457_o = ctrl[98:67]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:194:31  */
  assign n1459_o = 1'b1 ? n1457_o : rdata_gated;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:195:26  */
  assign n1460_o = ctrl[103]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:195:31  */
  assign n1462_o = 1'b1 ? n1460_o : ack_gated;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:196:26  */
  assign n1463_o = ctrl[104]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:196:31  */
  assign n1465_o = 1'b1 ? n1463_o : err_gated;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:140:5  */
  always @(posedge clk_i or posedge n1316_o)
    if (n1316_o)
      n1466_q <= n1411_o;
    else
      n1466_q <= n1409_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_xbus.vhd:129:5  */
  assign n1467_o = {n1465_o, n1462_o, n1459_o};
endmodule

module neorv32_bus_gateway_15_16384_8192_268435456_8192_8192_a510945699945b5d171ba29323e989d87bc97675
  (input  clk_i,
   input  rstn_i,
   input  [31:0] main_req_i_addr,
   input  [31:0] main_req_i_data,
   input  [3:0] main_req_i_ben,
   input  main_req_i_stb,
   input  main_req_i_rw,
   input  main_req_i_src,
   input  main_req_i_priv,
   input  main_req_i_rvso,
   input  main_req_i_fence,
   input  [31:0] imem_rsp_i_data,
   input  imem_rsp_i_ack,
   input  imem_rsp_i_err,
   input  [31:0] dmem_rsp_i_data,
   input  dmem_rsp_i_ack,
   input  dmem_rsp_i_err,
   input  [31:0] xip_rsp_i_data,
   input  xip_rsp_i_ack,
   input  xip_rsp_i_err,
   input  [31:0] boot_rsp_i_data,
   input  boot_rsp_i_ack,
   input  boot_rsp_i_err,
   input  [31:0] io_rsp_i_data,
   input  io_rsp_i_ack,
   input  io_rsp_i_err,
   input  [31:0] ext_rsp_i_data,
   input  ext_rsp_i_ack,
   input  ext_rsp_i_err,
   output [31:0] main_rsp_o_data,
   output main_rsp_o_ack,
   output main_rsp_o_err,
   output [31:0] imem_req_o_addr,
   output [31:0] imem_req_o_data,
   output [3:0] imem_req_o_ben,
   output imem_req_o_stb,
   output imem_req_o_rw,
   output imem_req_o_src,
   output imem_req_o_priv,
   output imem_req_o_rvso,
   output imem_req_o_fence,
   output [31:0] dmem_req_o_addr,
   output [31:0] dmem_req_o_data,
   output [3:0] dmem_req_o_ben,
   output dmem_req_o_stb,
   output dmem_req_o_rw,
   output dmem_req_o_src,
   output dmem_req_o_priv,
   output dmem_req_o_rvso,
   output dmem_req_o_fence,
   output [31:0] xip_req_o_addr,
   output [31:0] xip_req_o_data,
   output [3:0] xip_req_o_ben,
   output xip_req_o_stb,
   output xip_req_o_rw,
   output xip_req_o_src,
   output xip_req_o_priv,
   output xip_req_o_rvso,
   output xip_req_o_fence,
   output [31:0] boot_req_o_addr,
   output [31:0] boot_req_o_data,
   output [3:0] boot_req_o_ben,
   output boot_req_o_stb,
   output boot_req_o_rw,
   output boot_req_o_src,
   output boot_req_o_priv,
   output boot_req_o_rvso,
   output boot_req_o_fence,
   output [31:0] io_req_o_addr,
   output [31:0] io_req_o_data,
   output [3:0] io_req_o_ben,
   output io_req_o_stb,
   output io_req_o_rw,
   output io_req_o_src,
   output io_req_o_priv,
   output io_req_o_rvso,
   output io_req_o_fence,
   output [31:0] ext_req_o_addr,
   output [31:0] ext_req_o_data,
   output [3:0] ext_req_o_ben,
   output ext_req_o_stb,
   output ext_req_o_rw,
   output ext_req_o_src,
   output ext_req_o_priv,
   output ext_req_o_rvso,
   output ext_req_o_fence);
  wire [73:0] n1048_o;
  wire [31:0] n1050_o;
  wire n1051_o;
  wire n1052_o;
  wire [31:0] n1054_o;
  wire [31:0] n1055_o;
  wire [3:0] n1056_o;
  wire n1057_o;
  wire n1058_o;
  wire n1059_o;
  wire n1060_o;
  wire n1061_o;
  wire n1062_o;
  wire [33:0] n1063_o;
  wire [31:0] n1065_o;
  wire [31:0] n1066_o;
  wire [3:0] n1067_o;
  wire n1068_o;
  wire n1069_o;
  wire n1070_o;
  wire n1071_o;
  wire n1072_o;
  wire n1073_o;
  wire [33:0] n1074_o;
  wire [31:0] n1076_o;
  wire [31:0] n1077_o;
  wire [3:0] n1078_o;
  wire n1079_o;
  wire n1080_o;
  wire n1081_o;
  wire n1082_o;
  wire n1083_o;
  wire n1084_o;
  wire [33:0] n1085_o;
  wire [31:0] n1087_o;
  wire [31:0] n1088_o;
  wire [3:0] n1089_o;
  wire n1090_o;
  wire n1091_o;
  wire n1092_o;
  wire n1093_o;
  wire n1094_o;
  wire n1095_o;
  wire [33:0] n1096_o;
  wire [31:0] n1098_o;
  wire [31:0] n1099_o;
  wire [3:0] n1100_o;
  wire n1101_o;
  wire n1102_o;
  wire n1103_o;
  wire n1104_o;
  wire n1105_o;
  wire n1106_o;
  wire [33:0] n1107_o;
  wire [31:0] n1109_o;
  wire [31:0] n1110_o;
  wire [3:0] n1111_o;
  wire n1112_o;
  wire n1113_o;
  wire n1114_o;
  wire n1115_o;
  wire n1116_o;
  wire n1117_o;
  wire [33:0] n1118_o;
  wire [5:0] port_sel;
  wire [443:0] port_req;
  wire [203:0] port_rsp;
  wire [33:0] int_rsp;
  wire [7:0] keeper;
  wire n1126_o;
  wire n1135_o;
  wire n1144_o;
  wire n1153_o;
  wire [18:0] n1157_o;
  wire n1160_o;
  wire n1162_o;
  wire n1163_o;
  wire [4:0] n1166_o;
  wire n1168_o;
  wire n1170_o;
  wire n1171_o;
  wire [73:0] n1173_o;
  wire [73:0] n1174_o;
  wire [73:0] n1175_o;
  wire [73:0] n1176_o;
  wire [73:0] n1177_o;
  wire [73:0] n1178_o;
  wire n1181_o;
  wire n1182_o;
  wire n1183_o;
  wire [4:0] n1184_o;
  wire [67:0] n1185_o;
  wire n1186_o;
  wire n1187_o;
  wire n1188_o;
  wire [4:0] n1189_o;
  wire [67:0] n1190_o;
  localparam [33:0] n1194_o = 34'b0000000000000000000000000000000000;
  wire [31:0] n1195_o;
  wire [31:0] n1197_o;
  wire [31:0] n1198_o;
  localparam [33:0] n1199_o = 34'b0000000000000000000000000000000000;
  wire [1:0] n1200_o;
  wire [33:0] n1201_o;
  wire n1202_o;
  wire n1204_o;
  wire n1205_o;
  wire n1206_o;
  wire [33:0] n1207_o;
  wire n1208_o;
  wire n1210_o;
  wire n1211_o;
  wire [33:0] n1212_o;
  wire [31:0] n1213_o;
  wire [31:0] n1215_o;
  wire [31:0] n1216_o;
  wire [33:0] n1217_o;
  wire n1218_o;
  wire n1220_o;
  wire n1221_o;
  wire [33:0] n1222_o;
  wire n1223_o;
  wire n1225_o;
  wire n1226_o;
  wire [33:0] n1227_o;
  wire [31:0] n1230_o;
  wire n1231_o;
  wire n1232_o;
  wire n1234_o;
  wire n1241_o;
  wire n1242_o;
  wire n1243_o;
  wire n1244_o;
  wire n1245_o;
  wire n1247_o;
  wire [4:0] n1248_o;
  wire [4:0] n1250_o;
  wire n1251_o;
  wire n1259_o;
  wire n1261_o;
  wire n1263_o;
  wire n1264_o;
  wire n1265_o;
  wire n1266_o;
  wire n1267_o;
  wire n1268_o;
  wire n1269_o;
  wire n1270_o;
  wire n1271_o;
  wire n1272_o;
  wire n1273_o;
  wire n1274_o;
  wire n1275_o;
  wire n1278_o;
  wire n1280_o;
  wire n1281_o;
  wire n1282_o;
  wire n1283_o;
  wire [6:0] n1284_o;
  wire [5:0] n1285_o;
  wire [5:0] n1286_o;
  wire [5:0] n1287_o;
  wire n1288_o;
  wire n1289_o;
  wire [7:0] n1290_o;
  wire [7:0] n1292_o;
  wire [5:0] n1295_o;
  wire [443:0] n1296_o;
  wire [203:0] n1297_o;
  reg [7:0] n1298_q;
  wire [33:0] n1299_o;
  assign main_rsp_o_data = n1050_o; //(module output)
  assign main_rsp_o_ack = n1051_o; //(module output)
  assign main_rsp_o_err = n1052_o; //(module output)
  assign imem_req_o_addr = n1054_o; //(module output)
  assign imem_req_o_data = n1055_o; //(module output)
  assign imem_req_o_ben = n1056_o; //(module output)
  assign imem_req_o_stb = n1057_o; //(module output)
  assign imem_req_o_rw = n1058_o; //(module output)
  assign imem_req_o_src = n1059_o; //(module output)
  assign imem_req_o_priv = n1060_o; //(module output)
  assign imem_req_o_rvso = n1061_o; //(module output)
  assign imem_req_o_fence = n1062_o; //(module output)
  assign dmem_req_o_addr = n1065_o; //(module output)
  assign dmem_req_o_data = n1066_o; //(module output)
  assign dmem_req_o_ben = n1067_o; //(module output)
  assign dmem_req_o_stb = n1068_o; //(module output)
  assign dmem_req_o_rw = n1069_o; //(module output)
  assign dmem_req_o_src = n1070_o; //(module output)
  assign dmem_req_o_priv = n1071_o; //(module output)
  assign dmem_req_o_rvso = n1072_o; //(module output)
  assign dmem_req_o_fence = n1073_o; //(module output)
  assign xip_req_o_addr = n1076_o; //(module output)
  assign xip_req_o_data = n1077_o; //(module output)
  assign xip_req_o_ben = n1078_o; //(module output)
  assign xip_req_o_stb = n1079_o; //(module output)
  assign xip_req_o_rw = n1080_o; //(module output)
  assign xip_req_o_src = n1081_o; //(module output)
  assign xip_req_o_priv = n1082_o; //(module output)
  assign xip_req_o_rvso = n1083_o; //(module output)
  assign xip_req_o_fence = n1084_o; //(module output)
  assign boot_req_o_addr = n1087_o; //(module output)
  assign boot_req_o_data = n1088_o; //(module output)
  assign boot_req_o_ben = n1089_o; //(module output)
  assign boot_req_o_stb = n1090_o; //(module output)
  assign boot_req_o_rw = n1091_o; //(module output)
  assign boot_req_o_src = n1092_o; //(module output)
  assign boot_req_o_priv = n1093_o; //(module output)
  assign boot_req_o_rvso = n1094_o; //(module output)
  assign boot_req_o_fence = n1095_o; //(module output)
  assign io_req_o_addr = n1098_o; //(module output)
  assign io_req_o_data = n1099_o; //(module output)
  assign io_req_o_ben = n1100_o; //(module output)
  assign io_req_o_stb = n1101_o; //(module output)
  assign io_req_o_rw = n1102_o; //(module output)
  assign io_req_o_src = n1103_o; //(module output)
  assign io_req_o_priv = n1104_o; //(module output)
  assign io_req_o_rvso = n1105_o; //(module output)
  assign io_req_o_fence = n1106_o; //(module output)
  assign ext_req_o_addr = n1109_o; //(module output)
  assign ext_req_o_data = n1110_o; //(module output)
  assign ext_req_o_ben = n1111_o; //(module output)
  assign ext_req_o_stb = n1112_o; //(module output)
  assign ext_req_o_rw = n1113_o; //(module output)
  assign ext_req_o_src = n1114_o; //(module output)
  assign ext_req_o_priv = n1115_o; //(module output)
  assign ext_req_o_rvso = n1116_o; //(module output)
  assign ext_req_o_fence = n1117_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:55:5  */
  assign n1048_o = {main_req_i_fence, main_req_i_rvso, main_req_i_priv, main_req_i_src, main_req_i_rw, main_req_i_stb, main_req_i_ben, main_req_i_data, main_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:290:20  */
  assign n1050_o = n1299_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:94:3  */
  assign n1051_o = n1299_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1034:14  */
  assign n1052_o = n1299_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:451:13  */
  assign n1054_o = n1173_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:80:3  */
  assign n1055_o = n1173_o[63:32]; // extract
  assign n1056_o = n1173_o[67:64]; // extract
  assign n1057_o = n1173_o[68]; // extract
  assign n1058_o = n1173_o[69]; // extract
  assign n1059_o = n1173_o[70]; // extract
  assign n1060_o = n1173_o[71]; // extract
  assign n1061_o = n1173_o[72]; // extract
  assign n1062_o = n1173_o[73]; // extract
  assign n1063_o = {imem_rsp_i_err, imem_rsp_i_ack, imem_rsp_i_data};
  assign n1065_o = n1174_o[31:0]; // extract
  assign n1066_o = n1174_o[63:32]; // extract
  assign n1067_o = n1174_o[67:64]; // extract
  assign n1068_o = n1174_o[68]; // extract
  assign n1069_o = n1174_o[69]; // extract
  assign n1070_o = n1174_o[70]; // extract
  assign n1071_o = n1174_o[71]; // extract
  assign n1072_o = n1174_o[72]; // extract
  assign n1073_o = n1174_o[73]; // extract
  assign n1074_o = {dmem_rsp_i_err, dmem_rsp_i_ack, dmem_rsp_i_data};
  assign n1076_o = n1175_o[31:0]; // extract
  assign n1077_o = n1175_o[63:32]; // extract
  assign n1078_o = n1175_o[67:64]; // extract
  assign n1079_o = n1175_o[68]; // extract
  assign n1080_o = n1175_o[69]; // extract
  assign n1081_o = n1175_o[70]; // extract
  assign n1082_o = n1175_o[71]; // extract
  assign n1083_o = n1175_o[72]; // extract
  assign n1084_o = n1175_o[73]; // extract
  assign n1085_o = {xip_rsp_i_err, xip_rsp_i_ack, xip_rsp_i_data};
  assign n1087_o = n1176_o[31:0]; // extract
  assign n1088_o = n1176_o[63:32]; // extract
  assign n1089_o = n1176_o[67:64]; // extract
  assign n1090_o = n1176_o[68]; // extract
  assign n1091_o = n1176_o[69]; // extract
  assign n1092_o = n1176_o[70]; // extract
  assign n1093_o = n1176_o[71]; // extract
  assign n1094_o = n1176_o[72]; // extract
  assign n1095_o = n1176_o[73]; // extract
  assign n1096_o = {boot_rsp_i_err, boot_rsp_i_ack, boot_rsp_i_data};
  assign n1098_o = n1177_o[31:0]; // extract
  assign n1099_o = n1177_o[63:32]; // extract
  assign n1100_o = n1177_o[67:64]; // extract
  assign n1101_o = n1177_o[68]; // extract
  assign n1102_o = n1177_o[69]; // extract
  assign n1103_o = n1177_o[70]; // extract
  assign n1104_o = n1177_o[71]; // extract
  assign n1105_o = n1177_o[72]; // extract
  assign n1106_o = n1177_o[73]; // extract
  assign n1107_o = {io_rsp_i_err, io_rsp_i_ack, io_rsp_i_data};
  assign n1109_o = n1178_o[31:0]; // extract
  assign n1110_o = n1178_o[63:32]; // extract
  assign n1111_o = n1178_o[67:64]; // extract
  assign n1112_o = n1178_o[68]; // extract
  assign n1113_o = n1178_o[69]; // extract
  assign n1114_o = n1178_o[70]; // extract
  assign n1115_o = n1178_o[71]; // extract
  assign n1116_o = n1178_o[72]; // extract
  assign n1117_o = n1178_o[73]; // extract
  assign n1118_o = {ext_rsp_i_err, ext_rsp_i_ack, ext_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:274:10  */
  assign port_sel = n1295_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:283:10  */
  assign port_req = n1296_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:284:10  */
  assign port_rsp = n1297_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:287:10  */
  assign int_rsp = n1227_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:296:10  */
  assign keeper = n1298_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:302:22  */
  assign n1126_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:303:22  */
  assign n1135_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:304:22  */
  assign n1144_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:305:22  */
  assign n1153_o = 1'b0 ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:306:43  */
  assign n1157_o = n1048_o[31:13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:306:79  */
  assign n1160_o = n1157_o == 19'b1111111111111111111;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:306:127  */
  assign n1162_o = 1'b1 & n1160_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:306:22  */
  assign n1163_o = n1162_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:309:37  */
  assign n1166_o = port_sel[4:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:309:50  */
  assign n1168_o = n1166_o == 5'b00000;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:309:61  */
  assign n1170_o = 1'b1 & n1168_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:309:22  */
  assign n1171_o = n1170_o ? 1'b1 : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:314:25  */
  assign n1173_o = port_req[443:370]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:315:25  */
  assign n1174_o = port_req[369:296]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:316:25  */
  assign n1175_o = port_req[295:222]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:317:25  */
  assign n1176_o = port_req[221:148]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:318:25  */
  assign n1177_o = port_req[147:74]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:319:25  */
  assign n1178_o = port_req[73:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:328:39  */
  assign n1181_o = n1048_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:328:55  */
  assign n1182_o = port_sel[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:328:43  */
  assign n1183_o = n1181_o & n1182_o;
  assign n1184_o = n1048_o[73:69]; // extract
  assign n1185_o = n1048_o[67:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:328:39  */
  assign n1186_o = n1048_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:328:55  */
  assign n1187_o = port_sel[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:328:43  */
  assign n1188_o = n1186_o & n1187_o;
  assign n1189_o = n1048_o[73:69]; // extract
  assign n1190_o = n1048_o[67:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:340:29  */
  assign n1195_o = n1194_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:340:49  */
  assign n1197_o = port_rsp[65:34]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:340:34  */
  assign n1198_o = n1195_o | n1197_o;
  assign n1200_o = n1199_o[33:32]; // extract
  assign n1201_o = {n1200_o, n1198_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:341:29  */
  assign n1202_o = n1201_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:341:49  */
  assign n1204_o = port_rsp[66]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:341:34  */
  assign n1205_o = n1202_o | n1204_o;
  assign n1206_o = n1199_o[33]; // extract
  assign n1207_o = {n1206_o, n1205_o, n1198_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:342:29  */
  assign n1208_o = n1207_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:342:49  */
  assign n1210_o = port_rsp[67]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:342:34  */
  assign n1211_o = n1208_o | n1210_o;
  assign n1212_o = {n1211_o, n1205_o, n1198_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:340:29  */
  assign n1213_o = n1212_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:340:49  */
  assign n1215_o = port_rsp[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:340:34  */
  assign n1216_o = n1213_o | n1215_o;
  assign n1217_o = {n1211_o, n1205_o, n1216_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:341:29  */
  assign n1218_o = n1217_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:341:49  */
  assign n1220_o = port_rsp[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:341:34  */
  assign n1221_o = n1218_o | n1220_o;
  assign n1222_o = {n1211_o, n1221_o, n1216_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:342:29  */
  assign n1223_o = n1222_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:342:49  */
  assign n1225_o = port_rsp[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:342:34  */
  assign n1226_o = n1223_o | n1225_o;
  assign n1227_o = {n1226_o, n1221_o, n1216_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:349:30  */
  assign n1230_o = int_rsp[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:350:30  */
  assign n1231_o = int_rsp[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:351:29  */
  assign n1232_o = keeper[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:358:16  */
  assign n1234_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:365:30  */
  assign n1241_o = port_sel[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:365:45  */
  assign n1242_o = port_sel[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:365:34  */
  assign n1243_o = n1241_o | n1242_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:366:18  */
  assign n1244_o = keeper[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:366:23  */
  assign n1245_o = ~n1244_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:368:35  */
  assign n1247_o = n1048_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:370:57  */
  assign n1248_o = keeper[5:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:370:62  */
  assign n1250_o = n1248_o - 5'b00001;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:371:21  */
  assign n1251_o = int_rsp[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1259_o = keeper[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1261_o = 1'b0 | n1259_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1263_o = keeper[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1264_o = n1261_o | n1263_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1265_o = keeper[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1266_o = n1264_o | n1265_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1267_o = keeper[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1268_o = n1266_o | n1267_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:30  */
  assign n1269_o = keeper[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1026:22  */
  assign n1270_o = n1268_o | n1269_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:371:61  */
  assign n1271_o = ~n1270_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:371:80  */
  assign n1272_o = keeper[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:371:85  */
  assign n1273_o = ~n1272_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:371:68  */
  assign n1274_o = n1273_o & n1271_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:371:32  */
  assign n1275_o = n1251_o | n1274_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:374:24  */
  assign n1278_o = int_rsp[32]; // extract
  assign n1280_o = keeper[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:374:9  */
  assign n1281_o = n1278_o ? 1'b0 : n1280_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:371:9  */
  assign n1282_o = n1275_o ? 1'b0 : n1281_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:371:9  */
  assign n1283_o = n1275_o ? 1'b1 : 1'b0;
  assign n1284_o = {n1283_o, n1250_o, n1282_o};
  assign n1285_o = {5'b01111, n1247_o};
  assign n1286_o = n1284_o[5:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:366:7  */
  assign n1287_o = n1245_o ? n1285_o : n1286_o;
  assign n1288_o = n1284_o[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:366:7  */
  assign n1289_o = n1245_o ? 1'b0 : n1288_o;
  assign n1290_o = {n1243_o, n1289_o, n1287_o};
  assign n1292_o = {1'b0, 1'b0, 5'b00000, 1'b0};
  assign n1295_o = {n1171_o, n1163_o, n1153_o, n1144_o, n1135_o, n1126_o};
  assign n1296_o = {74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, 74'b00000000000000000000000000000000000000000000000000000000000000000000000000, n1184_o, n1183_o, n1185_o, n1189_o, n1188_o, n1190_o};
  assign n1297_o = {n1063_o, n1074_o, n1085_o, n1096_o, n1107_o, n1118_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:363:5  */
  always @(posedge clk_i or posedge n1234_o)
    if (n1234_o)
      n1298_q <= n1292_o;
    else
      n1298_q <= n1290_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:358:5  */
  assign n1299_o = {n1232_o, n1231_o, n1230_o};
endmodule

module neorv32_bus_switch_3f29546453678b855931c174a97d6c0894b8f546
  (input  clk_i,
   input  rstn_i,
   input  [31:0] a_req_i_addr,
   input  [31:0] a_req_i_data,
   input  [3:0] a_req_i_ben,
   input  a_req_i_stb,
   input  a_req_i_rw,
   input  a_req_i_src,
   input  a_req_i_priv,
   input  a_req_i_rvso,
   input  a_req_i_fence,
   input  [31:0] b_req_i_addr,
   input  [31:0] b_req_i_data,
   input  [3:0] b_req_i_ben,
   input  b_req_i_stb,
   input  b_req_i_rw,
   input  b_req_i_src,
   input  b_req_i_priv,
   input  b_req_i_rvso,
   input  b_req_i_fence,
   input  [31:0] x_rsp_i_data,
   input  x_rsp_i_ack,
   input  x_rsp_i_err,
   output [31:0] a_rsp_o_data,
   output a_rsp_o_ack,
   output a_rsp_o_err,
   output [31:0] b_rsp_o_data,
   output b_rsp_o_ack,
   output b_rsp_o_err,
   output [31:0] x_req_o_addr,
   output [31:0] x_req_o_data,
   output [3:0] x_req_o_ben,
   output x_req_o_stb,
   output x_req_o_rw,
   output x_req_o_src,
   output x_req_o_priv,
   output x_req_o_rvso,
   output x_req_o_fence);
  wire [73:0] n877_o;
  wire [31:0] n879_o;
  wire n880_o;
  wire n881_o;
  wire [73:0] n882_o;
  wire [31:0] n884_o;
  wire n885_o;
  wire n886_o;
  wire [31:0] n888_o;
  wire [31:0] n889_o;
  wire [3:0] n890_o;
  wire n891_o;
  wire n892_o;
  wire n893_o;
  wire n894_o;
  wire n895_o;
  wire n896_o;
  wire [33:0] n897_o;
  wire [7:0] arbiter;
  wire n899_o;
  wire [1:0] n904_o;
  wire n905_o;
  wire n906_o;
  wire n907_o;
  wire n908_o;
  wire n909_o;
  wire n910_o;
  wire n911_o;
  wire n912_o;
  wire n913_o;
  wire n914_o;
  wire n915_o;
  wire n916_o;
  wire [1:0] n917_o;
  wire [1:0] n922_o;
  wire [1:0] n927_o;
  wire [1:0] n930_o;
  wire n932_o;
  wire n933_o;
  wire n934_o;
  wire [1:0] n935_o;
  wire n937_o;
  wire n939_o;
  wire n940_o;
  wire n941_o;
  wire [1:0] n942_o;
  wire n944_o;
  wire n945_o;
  wire n946_o;
  wire n947_o;
  wire n951_o;
  wire n952_o;
  wire n953_o;
  wire [1:0] n957_o;
  wire [1:0] n958_o;
  wire [1:0] n959_o;
  wire [1:0] n960_o;
  wire [1:0] n961_o;
  wire [1:0] n962_o;
  wire [1:0] n963_o;
  wire [1:0] n964_o;
  reg [1:0] n965_o;
  wire n966_o;
  reg n967_o;
  wire n968_o;
  reg n969_o;
  wire [31:0] n971_o;
  wire n972_o;
  wire n973_o;
  wire [31:0] n974_o;
  wire [31:0] n975_o;
  wire n976_o;
  wire n977_o;
  wire n978_o;
  wire n979_o;
  wire n980_o;
  wire n981_o;
  wire n982_o;
  wire n983_o;
  wire n984_o;
  wire n985_o;
  wire n986_o;
  wire n987_o;
  wire n988_o;
  wire n989_o;
  wire n990_o;
  wire n991_o;
  wire n992_o;
  wire n993_o;
  wire n994_o;
  wire n995_o;
  wire n996_o;
  wire n997_o;
  wire n998_o;
  wire [31:0] n999_o;
  wire [31:0] n1001_o;
  wire [31:0] n1002_o;
  wire [31:0] n1004_o;
  wire [31:0] n1005_o;
  wire n1006_o;
  wire n1007_o;
  wire [31:0] n1008_o;
  wire [31:0] n1009_o;
  wire [3:0] n1010_o;
  wire [3:0] n1012_o;
  wire [3:0] n1013_o;
  wire [3:0] n1015_o;
  wire [3:0] n1016_o;
  wire n1017_o;
  wire n1018_o;
  wire [3:0] n1019_o;
  wire [3:0] n1020_o;
  wire n1021_o;
  wire [31:0] n1022_o;
  wire n1023_o;
  wire n1024_o;
  wire n1025_o;
  wire n1026_o;
  wire n1028_o;
  wire n1029_o;
  wire n1030_o;
  wire n1031_o;
  wire [31:0] n1033_o;
  wire n1034_o;
  wire n1035_o;
  wire n1036_o;
  wire n1038_o;
  wire n1039_o;
  wire n1040_o;
  reg [1:0] n1042_q;
  reg [1:0] n1043_q;
  wire [7:0] n1044_o;
  wire [33:0] n1045_o;
  wire [33:0] n1046_o;
  wire [73:0] n1047_o;
  assign a_rsp_o_data = n879_o; //(module output)
  assign a_rsp_o_ack = n880_o; //(module output)
  assign a_rsp_o_err = n881_o; //(module output)
  assign b_rsp_o_data = n884_o; //(module output)
  assign b_rsp_o_ack = n885_o; //(module output)
  assign b_rsp_o_err = n886_o; //(module output)
  assign x_req_o_addr = n888_o; //(module output)
  assign x_req_o_data = n889_o; //(module output)
  assign x_req_o_ben = n890_o; //(module output)
  assign x_req_o_stb = n891_o; //(module output)
  assign x_req_o_rw = n892_o; //(module output)
  assign x_req_o_src = n893_o; //(module output)
  assign x_req_o_priv = n894_o; //(module output)
  assign x_req_o_rvso = n895_o; //(module output)
  assign x_req_o_fence = n896_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:343:20  */
  assign n877_o = {a_req_i_fence, a_req_i_rvso, a_req_i_priv, a_req_i_src, a_req_i_rw, a_req_i_stb, a_req_i_ben, a_req_i_data, a_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:341:20  */
  assign n879_o = n1045_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:340:20  */
  assign n880_o = n1045_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:339:20  */
  assign n881_o = n1045_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:338:20  */
  assign n882_o = {b_req_i_fence, b_req_i_rvso, b_req_i_priv, b_req_i_src, b_req_i_rw, b_req_i_stb, b_req_i_ben, b_req_i_data, b_req_i_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:319:20  */
  assign n884_o = n1046_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:317:20  */
  assign n885_o = n1046_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:316:20  */
  assign n886_o = n1046_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:306:20  */
  assign n888_o = n1047_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:278:15  */
  assign n889_o = n1047_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:277:15  */
  assign n890_o = n1047_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:276:15  */
  assign n891_o = n1047_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:275:15  */
  assign n892_o = n1047_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:230:22  */
  assign n893_o = n1047_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:229:22  */
  assign n894_o = n1047_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:228:22  */
  assign n895_o = n1047_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:226:22  */
  assign n896_o = n1047_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:225:22  */
  assign n897_o = {x_rsp_i_err, x_rsp_i_ack, x_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:69:10  */
  assign arbiter = n1044_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:82:16  */
  assign n899_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:87:32  */
  assign n904_o = arbiter[3:2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:33  */
  assign n905_o = arbiter[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:50  */
  assign n906_o = n877_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:39  */
  assign n907_o = n905_o | n906_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:77  */
  assign n908_o = arbiter[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:60  */
  assign n909_o = ~n908_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:88:55  */
  assign n910_o = n907_o & n909_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:33  */
  assign n911_o = arbiter[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:50  */
  assign n912_o = n882_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:39  */
  assign n913_o = n911_o | n912_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:77  */
  assign n914_o = arbiter[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:60  */
  assign n915_o = ~n914_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:89:55  */
  assign n916_o = n913_o & n915_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:452:25  */
  assign n917_o = {n916_o, n910_o};
  assign n922_o = {1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:97:34  */
  assign n927_o = arbiter[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:102:18  */
  assign n930_o = arbiter[1:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:107:21  */
  assign n932_o = n897_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:107:44  */
  assign n933_o = n897_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:107:32  */
  assign n934_o = n932_o | n933_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:107:9  */
  assign n935_o = n934_o ? 2'b00 : n927_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:104:7  */
  assign n937_o = n930_o == 2'b01;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:114:21  */
  assign n939_o = n897_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:114:44  */
  assign n940_o = n897_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:114:32  */
  assign n941_o = n939_o | n940_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:114:9  */
  assign n942_o = n941_o ? 2'b00 : n927_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:111:7  */
  assign n944_o = n930_o == 2'b10;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:21  */
  assign n945_o = n877_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:44  */
  assign n946_o = arbiter[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:32  */
  assign n947_o = n945_o | n946_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:24  */
  assign n951_o = n882_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:47  */
  assign n952_o = arbiter[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:35  */
  assign n953_o = n951_o | n952_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:325:31  */
  assign n957_o = {1'b1, 1'b1};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:9  */
  assign n958_o = n953_o ? 2'b10 : n927_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:310:10  */
  assign n959_o = {1'b0, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:124:9  */
  assign n960_o = n953_o ? n957_o : n959_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:306:21  */
  assign n961_o = {1'b1, 1'b0};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:9  */
  assign n962_o = n947_o ? 2'b01 : n958_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:120:9  */
  assign n963_o = n947_o ? n961_o : n960_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:297:22  */
  assign n964_o = {n944_o, n937_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:102:5  */
  always @*
    case (n964_o)
      2'b10: n965_o = n942_o;
      2'b01: n965_o = n935_o;
      default: n965_o = n962_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:296:10  */
  assign n966_o = n963_o[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:102:5  */
  always @*
    case (n964_o)
      2'b10: n967_o = 1'b1;
      2'b01: n967_o = 1'b0;
      default: n967_o = n966_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:295:10  */
  assign n968_o = n963_o[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:102:5  */
  always @*
    case (n964_o)
      2'b10: n969_o = 1'b0;
      2'b01: n969_o = 1'b0;
      default: n969_o = n968_o;
    endcase
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:28  */
  assign n971_o = n877_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:47  */
  assign n972_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:51  */
  assign n973_o = ~n972_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:33  */
  assign n974_o = n973_o ? n971_o : n975_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:136:71  */
  assign n975_o = n882_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:28  */
  assign n976_o = n877_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:47  */
  assign n977_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:51  */
  assign n978_o = ~n977_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:33  */
  assign n979_o = n978_o ? n976_o : n980_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:137:71  */
  assign n980_o = n882_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:28  */
  assign n981_o = n877_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:47  */
  assign n982_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:51  */
  assign n983_o = ~n982_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:33  */
  assign n984_o = n983_o ? n981_o : n985_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:138:71  */
  assign n985_o = n882_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:28  */
  assign n986_o = n877_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:47  */
  assign n987_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:51  */
  assign n988_o = ~n987_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:33  */
  assign n989_o = n988_o ? n986_o : n990_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:139:71  */
  assign n990_o = n882_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:28  */
  assign n991_o = n877_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:47  */
  assign n992_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:51  */
  assign n993_o = ~n992_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:33  */
  assign n994_o = n993_o ? n991_o : n995_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:140:71  */
  assign n995_o = n882_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:141:28  */
  assign n996_o = n877_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:141:45  */
  assign n997_o = n882_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:141:34  */
  assign n998_o = n996_o | n997_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:143:28  */
  assign n999_o = n882_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:143:33  */
  assign n1001_o = 1'b0 ? n999_o : n1004_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:144:28  */
  assign n1002_o = n877_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:143:58  */
  assign n1004_o = 1'b1 ? n1002_o : n1008_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:145:28  */
  assign n1005_o = n877_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:145:47  */
  assign n1006_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:145:51  */
  assign n1007_o = ~n1006_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:144:58  */
  assign n1008_o = n1007_o ? n1005_o : n1009_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:145:71  */
  assign n1009_o = n882_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:147:28  */
  assign n1010_o = n882_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:147:32  */
  assign n1012_o = 1'b0 ? n1010_o : n1015_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:148:28  */
  assign n1013_o = n877_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:147:58  */
  assign n1015_o = 1'b1 ? n1013_o : n1019_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:149:28  */
  assign n1016_o = n877_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:149:46  */
  assign n1017_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:149:50  */
  assign n1018_o = ~n1017_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:148:58  */
  assign n1019_o = n1018_o ? n1016_o : n1020_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:149:71  */
  assign n1020_o = n882_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:151:28  */
  assign n1021_o = arbiter[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:156:27  */
  assign n1022_o = n897_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:157:27  */
  assign n1023_o = n897_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:157:45  */
  assign n1024_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:157:49  */
  assign n1025_o = ~n1024_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:157:31  */
  assign n1026_o = n1025_o ? n1023_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:158:27  */
  assign n1028_o = n897_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:158:45  */
  assign n1029_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:158:49  */
  assign n1030_o = ~n1029_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:158:31  */
  assign n1031_o = n1030_o ? n1028_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:160:27  */
  assign n1033_o = n897_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:161:27  */
  assign n1034_o = n897_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:161:45  */
  assign n1035_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:161:31  */
  assign n1036_o = n1035_o ? n1034_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:162:27  */
  assign n1038_o = n897_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:162:45  */
  assign n1039_o = arbiter[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:162:31  */
  assign n1040_o = n1039_o ? n1038_o : 1'b0;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:86:5  */
  always @(posedge clk_i or posedge n899_o)
    if (n899_o)
      n1042_q <= n922_o;
    else
      n1042_q <= n917_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:86:5  */
  always @(posedge clk_i or posedge n899_o)
    if (n899_o)
      n1043_q <= 2'b00;
    else
      n1043_q <= n904_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:82:5  */
  assign n1044_o = {n969_o, n967_o, n1042_q, n965_o, n1043_q};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_intercon.vhd:82:5  */
  assign n1045_o = {n1031_o, n1026_o, n1022_o};
  assign n1046_o = {n1040_o, n1036_o, n1033_o};
  assign n1047_o = {n998_o, n979_o, n984_o, n989_o, n994_o, n1021_o, n1012_o, n1001_o, n974_o};
endmodule

module neorv32_cpu_0_4_0_64_16973a3472ca3522cdc18159c73abb10ac4c9817
  (input  clk_i,
   input  clk_aux_i,
   input  rstn_i,
   input  msi_i,
   input  mei_i,
   input  mti_i,
   input  [15:0] firq_i,
   input  dbi_i,
   input  [31:0] ibus_rsp_i_data,
   input  ibus_rsp_i_ack,
   input  ibus_rsp_i_err,
   input  [31:0] dbus_rsp_i_data,
   input  dbus_rsp_i_ack,
   input  dbus_rsp_i_err,
   output sleep_o,
   output debug_o,
   output [31:0] ibus_req_o_addr,
   output [31:0] ibus_req_o_data,
   output [3:0] ibus_req_o_ben,
   output ibus_req_o_stb,
   output ibus_req_o_rw,
   output ibus_req_o_src,
   output ibus_req_o_priv,
   output ibus_req_o_rvso,
   output ibus_req_o_fence,
   output [31:0] dbus_req_o_addr,
   output [31:0] dbus_req_o_data,
   output [3:0] dbus_req_o_ben,
   output dbus_req_o_stb,
   output dbus_req_o_rw,
   output dbus_req_o_src,
   output dbus_req_o_priv,
   output dbus_req_o_rvso,
   output dbus_req_o_fence);
  wire [31:0] n722_o;
  wire [31:0] n723_o;
  wire [3:0] n724_o;
  wire n725_o;
  wire n726_o;
  wire n727_o;
  wire n728_o;
  wire n729_o;
  wire n730_o;
  wire [33:0] n731_o;
  wire [31:0] n733_o;
  wire [31:0] n734_o;
  wire [3:0] n735_o;
  wire n736_o;
  wire n737_o;
  wire n738_o;
  wire n739_o;
  wire n740_o;
  wire n741_o;
  wire [33:0] n742_o;
  wire xcsr_we;
  wire [11:0] xcsr_addr;
  wire [31:0] xcsr_wdata;
  wire [31:0] xcsr_rdata_pmp;
  wire [31:0] xcsr_rdata_alu;
  wire [31:0] xcsr_rdata_res;
  wire [66:0] ctrl;
  wire [31:0] imm;
  wire [31:0] rs1;
  wire [31:0] rs2;
  wire [31:0] rs3;
  wire [31:0] rs4;
  wire [31:0] alu_res;
  wire [31:0] alu_add;
  wire [1:0] alu_cmp;
  wire [31:0] mem_rdata;
  wire cp_done;
  wire lsu_wait;
  wire [31:0] csr_rdata;
  wire [31:0] mar;
  wire ma_load;
  wire ma_store;
  wire be_load;
  wire be_store;
  wire [31:0] curr_pc;
  wire [31:0] link_pc;
  wire pmp_ex_fault;
  wire pmp_rw_fault;
  wire neorv32_cpu_control_inst_ctrl_o_rf_wb_en;
  wire [4:0] neorv32_cpu_control_inst_ctrl_o_rf_rs1;
  wire [4:0] neorv32_cpu_control_inst_ctrl_o_rf_rs2;
  wire [4:0] neorv32_cpu_control_inst_ctrl_o_rf_rs3;
  wire [4:0] neorv32_cpu_control_inst_ctrl_o_rf_rd;
  wire [1:0] neorv32_cpu_control_inst_ctrl_o_rf_mux;
  wire neorv32_cpu_control_inst_ctrl_o_rf_zero_we;
  wire [2:0] neorv32_cpu_control_inst_ctrl_o_alu_op;
  wire neorv32_cpu_control_inst_ctrl_o_alu_opa_mux;
  wire neorv32_cpu_control_inst_ctrl_o_alu_opb_mux;
  wire neorv32_cpu_control_inst_ctrl_o_alu_unsigned;
  wire [5:0] neorv32_cpu_control_inst_ctrl_o_alu_cp_trig;
  wire neorv32_cpu_control_inst_ctrl_o_lsu_req;
  wire neorv32_cpu_control_inst_ctrl_o_lsu_rw;
  wire neorv32_cpu_control_inst_ctrl_o_lsu_mo_we;
  wire neorv32_cpu_control_inst_ctrl_o_lsu_fence;
  wire neorv32_cpu_control_inst_ctrl_o_lsu_priv;
  wire [2:0] neorv32_cpu_control_inst_ctrl_o_ir_funct3;
  wire [11:0] neorv32_cpu_control_inst_ctrl_o_ir_funct12;
  wire [6:0] neorv32_cpu_control_inst_ctrl_o_ir_opcode;
  wire neorv32_cpu_control_inst_ctrl_o_cpu_priv;
  wire neorv32_cpu_control_inst_ctrl_o_cpu_sleep;
  wire neorv32_cpu_control_inst_ctrl_o_cpu_trap;
  wire neorv32_cpu_control_inst_ctrl_o_cpu_debug;
  wire [31:0] neorv32_cpu_control_inst_bus_req_o_addr;
  wire [31:0] neorv32_cpu_control_inst_bus_req_o_data;
  wire [3:0] neorv32_cpu_control_inst_bus_req_o_ben;
  wire neorv32_cpu_control_inst_bus_req_o_stb;
  wire neorv32_cpu_control_inst_bus_req_o_rw;
  wire neorv32_cpu_control_inst_bus_req_o_src;
  wire neorv32_cpu_control_inst_bus_req_o_priv;
  wire neorv32_cpu_control_inst_bus_req_o_rvso;
  wire neorv32_cpu_control_inst_bus_req_o_fence;
  wire [31:0] neorv32_cpu_control_inst_imm_o;
  wire [31:0] neorv32_cpu_control_inst_fetch_pc_o;
  wire [31:0] neorv32_cpu_control_inst_curr_pc_o;
  wire [31:0] neorv32_cpu_control_inst_link_pc_o;
  wire [31:0] neorv32_cpu_control_inst_csr_rdata_o;
  wire neorv32_cpu_control_inst_xcsr_we_o;
  wire [11:0] neorv32_cpu_control_inst_xcsr_addr_o;
  wire [31:0] neorv32_cpu_control_inst_xcsr_wdata_o;
  wire [66:0] n763_o;
  wire [73:0] n765_o;
  wire [31:0] n767_o;
  wire n768_o;
  wire n769_o;
  wire [31:0] n778_o;
  wire n779_o;
  wire n780_o;
  wire [31:0] neorv32_cpu_regfile_inst_rs1_o;
  wire [31:0] neorv32_cpu_regfile_inst_rs2_o;
  wire [31:0] neorv32_cpu_regfile_inst_rs3_o;
  wire [31:0] neorv32_cpu_regfile_inst_rs4_o;
  wire n781_o;
  wire [4:0] n782_o;
  wire [4:0] n783_o;
  wire [4:0] n784_o;
  wire [4:0] n785_o;
  wire [1:0] n786_o;
  wire n787_o;
  wire [2:0] n788_o;
  wire n789_o;
  wire n790_o;
  wire n791_o;
  wire [5:0] n792_o;
  wire n793_o;
  wire n794_o;
  wire n795_o;
  wire n796_o;
  wire n797_o;
  wire [2:0] n798_o;
  wire [11:0] n799_o;
  wire [6:0] n800_o;
  wire n801_o;
  wire n802_o;
  wire n803_o;
  wire n804_o;
  wire [31:0] neorv32_cpu_alu_inst_csr_rdata_o;
  wire [1:0] neorv32_cpu_alu_inst_cmp_o;
  wire [31:0] neorv32_cpu_alu_inst_res_o;
  wire [31:0] neorv32_cpu_alu_inst_add_o;
  wire neorv32_cpu_alu_inst_cp_done_o;
  wire n809_o;
  wire [4:0] n810_o;
  wire [4:0] n811_o;
  wire [4:0] n812_o;
  wire [4:0] n813_o;
  wire [1:0] n814_o;
  wire n815_o;
  wire [2:0] n816_o;
  wire n817_o;
  wire n818_o;
  wire n819_o;
  wire [5:0] n820_o;
  wire n821_o;
  wire n822_o;
  wire n823_o;
  wire n824_o;
  wire n825_o;
  wire [2:0] n826_o;
  wire [11:0] n827_o;
  wire [6:0] n828_o;
  wire n829_o;
  wire n830_o;
  wire n831_o;
  wire n832_o;
  wire [31:0] neorv32_cpu_lsu_inst_rdata_o;
  wire [31:0] neorv32_cpu_lsu_inst_mar_o;
  wire neorv32_cpu_lsu_inst_wait_o;
  wire neorv32_cpu_lsu_inst_ma_load_o;
  wire neorv32_cpu_lsu_inst_ma_store_o;
  wire neorv32_cpu_lsu_inst_be_load_o;
  wire neorv32_cpu_lsu_inst_be_store_o;
  wire [31:0] neorv32_cpu_lsu_inst_bus_req_o_addr;
  wire [31:0] neorv32_cpu_lsu_inst_bus_req_o_data;
  wire [3:0] neorv32_cpu_lsu_inst_bus_req_o_ben;
  wire neorv32_cpu_lsu_inst_bus_req_o_stb;
  wire neorv32_cpu_lsu_inst_bus_req_o_rw;
  wire neorv32_cpu_lsu_inst_bus_req_o_src;
  wire neorv32_cpu_lsu_inst_bus_req_o_priv;
  wire neorv32_cpu_lsu_inst_bus_req_o_rvso;
  wire neorv32_cpu_lsu_inst_bus_req_o_fence;
  wire n838_o;
  wire [4:0] n839_o;
  wire [4:0] n840_o;
  wire [4:0] n841_o;
  wire [4:0] n842_o;
  wire [1:0] n843_o;
  wire n844_o;
  wire [2:0] n845_o;
  wire n846_o;
  wire n847_o;
  wire n848_o;
  wire [5:0] n849_o;
  wire n850_o;
  wire n851_o;
  wire n852_o;
  wire n853_o;
  wire n854_o;
  wire [2:0] n855_o;
  wire [11:0] n856_o;
  wire [6:0] n857_o;
  wire n858_o;
  wire n859_o;
  wire n860_o;
  wire n861_o;
  wire [73:0] n869_o;
  wire [31:0] n871_o;
  wire n872_o;
  wire n873_o;
  assign sleep_o = n779_o; //(module output)
  assign debug_o = n780_o; //(module output)
  assign ibus_req_o_addr = n722_o; //(module output)
  assign ibus_req_o_data = n723_o; //(module output)
  assign ibus_req_o_ben = n724_o; //(module output)
  assign ibus_req_o_stb = n725_o; //(module output)
  assign ibus_req_o_rw = n726_o; //(module output)
  assign ibus_req_o_src = n727_o; //(module output)
  assign ibus_req_o_priv = n728_o; //(module output)
  assign ibus_req_o_rvso = n729_o; //(module output)
  assign ibus_req_o_fence = n730_o; //(module output)
  assign dbus_req_o_addr = n733_o; //(module output)
  assign dbus_req_o_data = n734_o; //(module output)
  assign dbus_req_o_ben = n735_o; //(module output)
  assign dbus_req_o_stb = n736_o; //(module output)
  assign dbus_req_o_rw = n737_o; //(module output)
  assign dbus_req_o_src = n738_o; //(module output)
  assign dbus_req_o_priv = n739_o; //(module output)
  assign dbus_req_o_rvso = n740_o; //(module output)
  assign dbus_req_o_fence = n741_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1076:23  */
  assign n722_o = n765_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1075:23  */
  assign n723_o = n765_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1074:23  */
  assign n724_o = n765_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1073:23  */
  assign n725_o = n765_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1072:23  */
  assign n726_o = n765_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1071:23  */
  assign n727_o = n765_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1070:23  */
  assign n728_o = n765_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1069:23  */
  assign n729_o = n765_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1068:23  */
  assign n730_o = n765_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1067:23  */
  assign n731_o = {ibus_rsp_i_err, ibus_rsp_i_ack, ibus_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1065:23  */
  assign n733_o = n869_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1064:23  */
  assign n734_o = n869_o[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1063:23  */
  assign n735_o = n869_o[67:64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1062:23  */
  assign n736_o = n869_o[68]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1061:23  */
  assign n737_o = n869_o[69]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1060:23  */
  assign n738_o = n869_o[70]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1059:23  */
  assign n739_o = n869_o[71]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1058:23  */
  assign n740_o = n869_o[72]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1057:23  */
  assign n741_o = n869_o[73]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1056:23  */
  assign n742_o = {dbus_rsp_i_err, dbus_rsp_i_ack, dbus_rsp_i_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:107:10  */
  assign xcsr_we = neorv32_cpu_control_inst_xcsr_we_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:108:10  */
  assign xcsr_addr = neorv32_cpu_control_inst_xcsr_addr_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:109:10  */
  assign xcsr_wdata = neorv32_cpu_control_inst_xcsr_wdata_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:110:10  */
  assign xcsr_rdata_pmp = 32'b00000000000000000000000000000000; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:111:10  */
  assign xcsr_rdata_alu = neorv32_cpu_alu_inst_csr_rdata_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:112:10  */
  assign xcsr_rdata_res = n778_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:115:10  */
  assign ctrl = n763_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:116:10  */
  assign imm = neorv32_cpu_control_inst_imm_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:117:10  */
  assign rs1 = neorv32_cpu_regfile_inst_rs1_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:117:15  */
  assign rs2 = neorv32_cpu_regfile_inst_rs2_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:118:10  */
  assign rs3 = neorv32_cpu_regfile_inst_rs3_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:118:15  */
  assign rs4 = neorv32_cpu_regfile_inst_rs4_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:119:10  */
  assign alu_res = neorv32_cpu_alu_inst_res_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:120:10  */
  assign alu_add = neorv32_cpu_alu_inst_add_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:121:10  */
  assign alu_cmp = neorv32_cpu_alu_inst_cmp_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:122:10  */
  assign mem_rdata = neorv32_cpu_lsu_inst_rdata_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:123:10  */
  assign cp_done = neorv32_cpu_alu_inst_cp_done_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:124:10  */
  assign lsu_wait = neorv32_cpu_lsu_inst_wait_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:125:10  */
  assign csr_rdata = neorv32_cpu_control_inst_csr_rdata_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:126:10  */
  assign mar = neorv32_cpu_lsu_inst_mar_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:127:10  */
  assign ma_load = neorv32_cpu_lsu_inst_ma_load_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:128:10  */
  assign ma_store = neorv32_cpu_lsu_inst_ma_store_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:129:10  */
  assign be_load = neorv32_cpu_lsu_inst_be_load_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:130:10  */
  assign be_store = neorv32_cpu_lsu_inst_be_store_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:132:10  */
  assign curr_pc = neorv32_cpu_control_inst_curr_pc_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:133:10  */
  assign link_pc = neorv32_cpu_control_inst_link_pc_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:134:10  */
  assign pmp_ex_fault = 1'b0; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:135:10  */
  assign pmp_rw_fault = 1'b0; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:175:3  */
  neorv32_cpu_control_0_64_87d7d7036038d959ad02bd289905a845d3f42491 neorv32_cpu_control_inst (
    .clk_i(clk_i),
    .clk_aux_i(clk_aux_i),
    .rstn_i(rstn_i),
    .i_pmp_fault_i(pmp_ex_fault),
    .bus_rsp_i_data(n767_o),
    .bus_rsp_i_ack(n768_o),
    .bus_rsp_i_err(n769_o),
    .alu_cp_done_i(cp_done),
    .cmp_i(alu_cmp),
    .alu_add_i(alu_add),
    .rs1_i(rs1),
    .xcsr_rdata_i(xcsr_rdata_res),
    .db_halt_req_i(dbi_i),
    .msi_i(msi_i),
    .mei_i(mei_i),
    .mti_i(mti_i),
    .firq_i(firq_i),
    .lsu_wait_i(lsu_wait),
    .mar_i(mar),
    .ma_load_i(ma_load),
    .ma_store_i(ma_store),
    .be_load_i(be_load),
    .be_store_i(be_store),
    .ctrl_o_rf_wb_en(neorv32_cpu_control_inst_ctrl_o_rf_wb_en),
    .ctrl_o_rf_rs1(neorv32_cpu_control_inst_ctrl_o_rf_rs1),
    .ctrl_o_rf_rs2(neorv32_cpu_control_inst_ctrl_o_rf_rs2),
    .ctrl_o_rf_rs3(neorv32_cpu_control_inst_ctrl_o_rf_rs3),
    .ctrl_o_rf_rd(neorv32_cpu_control_inst_ctrl_o_rf_rd),
    .ctrl_o_rf_mux(neorv32_cpu_control_inst_ctrl_o_rf_mux),
    .ctrl_o_rf_zero_we(neorv32_cpu_control_inst_ctrl_o_rf_zero_we),
    .ctrl_o_alu_op(neorv32_cpu_control_inst_ctrl_o_alu_op),
    .ctrl_o_alu_opa_mux(neorv32_cpu_control_inst_ctrl_o_alu_opa_mux),
    .ctrl_o_alu_opb_mux(neorv32_cpu_control_inst_ctrl_o_alu_opb_mux),
    .ctrl_o_alu_unsigned(neorv32_cpu_control_inst_ctrl_o_alu_unsigned),
    .ctrl_o_alu_cp_trig(neorv32_cpu_control_inst_ctrl_o_alu_cp_trig),
    .ctrl_o_lsu_req(neorv32_cpu_control_inst_ctrl_o_lsu_req),
    .ctrl_o_lsu_rw(neorv32_cpu_control_inst_ctrl_o_lsu_rw),
    .ctrl_o_lsu_mo_we(neorv32_cpu_control_inst_ctrl_o_lsu_mo_we),
    .ctrl_o_lsu_fence(neorv32_cpu_control_inst_ctrl_o_lsu_fence),
    .ctrl_o_lsu_priv(neorv32_cpu_control_inst_ctrl_o_lsu_priv),
    .ctrl_o_ir_funct3(neorv32_cpu_control_inst_ctrl_o_ir_funct3),
    .ctrl_o_ir_funct12(neorv32_cpu_control_inst_ctrl_o_ir_funct12),
    .ctrl_o_ir_opcode(neorv32_cpu_control_inst_ctrl_o_ir_opcode),
    .ctrl_o_cpu_priv(neorv32_cpu_control_inst_ctrl_o_cpu_priv),
    .ctrl_o_cpu_sleep(neorv32_cpu_control_inst_ctrl_o_cpu_sleep),
    .ctrl_o_cpu_trap(neorv32_cpu_control_inst_ctrl_o_cpu_trap),
    .ctrl_o_cpu_debug(neorv32_cpu_control_inst_ctrl_o_cpu_debug),
    .bus_req_o_addr(neorv32_cpu_control_inst_bus_req_o_addr),
    .bus_req_o_data(neorv32_cpu_control_inst_bus_req_o_data),
    .bus_req_o_ben(neorv32_cpu_control_inst_bus_req_o_ben),
    .bus_req_o_stb(neorv32_cpu_control_inst_bus_req_o_stb),
    .bus_req_o_rw(neorv32_cpu_control_inst_bus_req_o_rw),
    .bus_req_o_src(neorv32_cpu_control_inst_bus_req_o_src),
    .bus_req_o_priv(neorv32_cpu_control_inst_bus_req_o_priv),
    .bus_req_o_rvso(neorv32_cpu_control_inst_bus_req_o_rvso),
    .bus_req_o_fence(neorv32_cpu_control_inst_bus_req_o_fence),
    .imm_o(neorv32_cpu_control_inst_imm_o),
    .fetch_pc_o(),
    .curr_pc_o(neorv32_cpu_control_inst_curr_pc_o),
    .link_pc_o(neorv32_cpu_control_inst_link_pc_o),
    .csr_rdata_o(neorv32_cpu_control_inst_csr_rdata_o),
    .xcsr_we_o(neorv32_cpu_control_inst_xcsr_we_o),
    .xcsr_addr_o(neorv32_cpu_control_inst_xcsr_addr_o),
    .xcsr_wdata_o(neorv32_cpu_control_inst_xcsr_wdata_o));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:212:5  */
  assign n763_o = {neorv32_cpu_control_inst_ctrl_o_cpu_debug, neorv32_cpu_control_inst_ctrl_o_cpu_trap, neorv32_cpu_control_inst_ctrl_o_cpu_sleep, neorv32_cpu_control_inst_ctrl_o_cpu_priv, neorv32_cpu_control_inst_ctrl_o_ir_opcode, neorv32_cpu_control_inst_ctrl_o_ir_funct12, neorv32_cpu_control_inst_ctrl_o_ir_funct3, neorv32_cpu_control_inst_ctrl_o_lsu_priv, neorv32_cpu_control_inst_ctrl_o_lsu_fence, neorv32_cpu_control_inst_ctrl_o_lsu_mo_we, neorv32_cpu_control_inst_ctrl_o_lsu_rw, neorv32_cpu_control_inst_ctrl_o_lsu_req, neorv32_cpu_control_inst_ctrl_o_alu_cp_trig, neorv32_cpu_control_inst_ctrl_o_alu_unsigned, neorv32_cpu_control_inst_ctrl_o_alu_opb_mux, neorv32_cpu_control_inst_ctrl_o_alu_opa_mux, neorv32_cpu_control_inst_ctrl_o_alu_op, neorv32_cpu_control_inst_ctrl_o_rf_zero_we, neorv32_cpu_control_inst_ctrl_o_rf_mux, neorv32_cpu_control_inst_ctrl_o_rf_rd, neorv32_cpu_control_inst_ctrl_o_rf_rs3, neorv32_cpu_control_inst_ctrl_o_rf_rs2, neorv32_cpu_control_inst_ctrl_o_rf_rs1, neorv32_cpu_control_inst_ctrl_o_rf_wb_en};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:206:5  */
  assign n765_o = {neorv32_cpu_control_inst_bus_req_o_fence, neorv32_cpu_control_inst_bus_req_o_rvso, neorv32_cpu_control_inst_bus_req_o_priv, neorv32_cpu_control_inst_bus_req_o_src, neorv32_cpu_control_inst_bus_req_o_rw, neorv32_cpu_control_inst_bus_req_o_stb, neorv32_cpu_control_inst_bus_req_o_ben, neorv32_cpu_control_inst_bus_req_o_data, neorv32_cpu_control_inst_bus_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:199:5  */
  assign n767_o = n731_o[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:197:5  */
  assign n768_o = n731_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:196:5  */
  assign n769_o = n731_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:248:36  */
  assign n778_o = xcsr_rdata_pmp | xcsr_rdata_alu;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:251:19  */
  assign n779_o = ctrl[64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:252:19  */
  assign n780_o = ctrl[66]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:257:3  */
  neorv32_cpu_regfile_9069ca78e7450a285173431b3e52c5c25299e473 neorv32_cpu_regfile_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n781_o),
    .ctrl_i_rf_rs1(n782_o),
    .ctrl_i_rf_rs2(n783_o),
    .ctrl_i_rf_rs3(n784_o),
    .ctrl_i_rf_rd(n785_o),
    .ctrl_i_rf_mux(n786_o),
    .ctrl_i_rf_zero_we(n787_o),
    .ctrl_i_alu_op(n788_o),
    .ctrl_i_alu_opa_mux(n789_o),
    .ctrl_i_alu_opb_mux(n790_o),
    .ctrl_i_alu_unsigned(n791_o),
    .ctrl_i_alu_cp_trig(n792_o),
    .ctrl_i_lsu_req(n793_o),
    .ctrl_i_lsu_rw(n794_o),
    .ctrl_i_lsu_mo_we(n795_o),
    .ctrl_i_lsu_fence(n796_o),
    .ctrl_i_lsu_priv(n797_o),
    .ctrl_i_ir_funct3(n798_o),
    .ctrl_i_ir_funct12(n799_o),
    .ctrl_i_ir_opcode(n800_o),
    .ctrl_i_cpu_priv(n801_o),
    .ctrl_i_cpu_sleep(n802_o),
    .ctrl_i_cpu_trap(n803_o),
    .ctrl_i_cpu_debug(n804_o),
    .alu_i(alu_res),
    .mem_i(mem_rdata),
    .csr_i(csr_rdata),
    .ret_i(link_pc),
    .rs1_o(neorv32_cpu_regfile_inst_rs1_o),
    .rs2_o(neorv32_cpu_regfile_inst_rs2_o),
    .rs3_o(neorv32_cpu_regfile_inst_rs3_o),
    .rs4_o(neorv32_cpu_regfile_inst_rs4_o));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:425:7  */
  assign n781_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:425:7  */
  assign n782_o = ctrl[5:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:425:7  */
  assign n783_o = ctrl[10:6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:449:7  */
  assign n784_o = ctrl[15:11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:465:7  */
  assign n785_o = ctrl[20:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:465:7  */
  assign n786_o = ctrl[22:21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:469:7  */
  assign n787_o = ctrl[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:465:7  */
  assign n788_o = ctrl[26:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:469:7  */
  assign n789_o = ctrl[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:469:7  */
  assign n790_o = ctrl[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:451:7  */
  assign n791_o = ctrl[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:430:7  */
  assign n792_o = ctrl[35:30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:430:7  */
  assign n793_o = ctrl[36]; // extract
  assign n794_o = ctrl[37]; // extract
  assign n795_o = ctrl[38]; // extract
  assign n796_o = ctrl[39]; // extract
  assign n797_o = ctrl[40]; // extract
  assign n798_o = ctrl[43:41]; // extract
  assign n799_o = ctrl[55:44]; // extract
  assign n800_o = ctrl[62:56]; // extract
  assign n801_o = ctrl[63]; // extract
  assign n802_o = ctrl[64]; // extract
  assign n803_o = ctrl[65]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1210:7  */
  assign n804_o = ctrl[66]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:284:3  */
  neorv32_cpu_alu_1db721083c34eba714927c673b29edb8e81e05fb neorv32_cpu_alu_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n809_o),
    .ctrl_i_rf_rs1(n810_o),
    .ctrl_i_rf_rs2(n811_o),
    .ctrl_i_rf_rs3(n812_o),
    .ctrl_i_rf_rd(n813_o),
    .ctrl_i_rf_mux(n814_o),
    .ctrl_i_rf_zero_we(n815_o),
    .ctrl_i_alu_op(n816_o),
    .ctrl_i_alu_opa_mux(n817_o),
    .ctrl_i_alu_opb_mux(n818_o),
    .ctrl_i_alu_unsigned(n819_o),
    .ctrl_i_alu_cp_trig(n820_o),
    .ctrl_i_lsu_req(n821_o),
    .ctrl_i_lsu_rw(n822_o),
    .ctrl_i_lsu_mo_we(n823_o),
    .ctrl_i_lsu_fence(n824_o),
    .ctrl_i_lsu_priv(n825_o),
    .ctrl_i_ir_funct3(n826_o),
    .ctrl_i_ir_funct12(n827_o),
    .ctrl_i_ir_opcode(n828_o),
    .ctrl_i_cpu_priv(n829_o),
    .ctrl_i_cpu_sleep(n830_o),
    .ctrl_i_cpu_trap(n831_o),
    .ctrl_i_cpu_debug(n832_o),
    .csr_we_i(xcsr_we),
    .csr_addr_i(xcsr_addr),
    .csr_wdata_i(xcsr_wdata),
    .rs1_i(rs1),
    .rs2_i(rs2),
    .rs3_i(rs3),
    .rs4_i(rs4),
    .pc_i(curr_pc),
    .imm_i(imm),
    .csr_rdata_o(neorv32_cpu_alu_inst_csr_rdata_o),
    .cmp_o(neorv32_cpu_alu_inst_cmp_o),
    .res_o(neorv32_cpu_alu_inst_res_o),
    .add_o(neorv32_cpu_alu_inst_add_o),
    .cp_done_o(neorv32_cpu_alu_inst_cp_done_o));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:801:19  */
  assign n809_o = ctrl[0]; // extract
  assign n810_o = ctrl[5:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:799:19  */
  assign n811_o = ctrl[10:6]; // extract
  assign n812_o = ctrl[15:11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:797:19  */
  assign n813_o = ctrl[20:16]; // extract
  assign n814_o = ctrl[22:21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:568:21  */
  assign n815_o = ctrl[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:567:21  */
  assign n816_o = ctrl[26:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:493:54  */
  assign n817_o = ctrl[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:493:62  */
  assign n818_o = ctrl[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:493:35  */
  assign n819_o = ctrl[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:493:43  */
  assign n820_o = ctrl[35:30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:492:93  */
  assign n821_o = ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:493:24  */
  assign n822_o = ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:492:73  */
  assign n823_o = ctrl[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:492:81  */
  assign n824_o = ctrl[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:492:54  */
  assign n825_o = ctrl[40]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:492:62  */
  assign n826_o = ctrl[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:492:35  */
  assign n827_o = ctrl[55:44]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:492:43  */
  assign n828_o = ctrl[62:56]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:491:93  */
  assign n829_o = ctrl[63]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:492:24  */
  assign n830_o = ctrl[64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:491:73  */
  assign n831_o = ctrl[65]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:491:81  */
  assign n832_o = ctrl[66]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_cpu.vhd:325:3  */
  neorv32_cpu_lsu_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_cpu_lsu_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .ctrl_i_rf_wb_en(n838_o),
    .ctrl_i_rf_rs1(n839_o),
    .ctrl_i_rf_rs2(n840_o),
    .ctrl_i_rf_rs3(n841_o),
    .ctrl_i_rf_rd(n842_o),
    .ctrl_i_rf_mux(n843_o),
    .ctrl_i_rf_zero_we(n844_o),
    .ctrl_i_alu_op(n845_o),
    .ctrl_i_alu_opa_mux(n846_o),
    .ctrl_i_alu_opb_mux(n847_o),
    .ctrl_i_alu_unsigned(n848_o),
    .ctrl_i_alu_cp_trig(n849_o),
    .ctrl_i_lsu_req(n850_o),
    .ctrl_i_lsu_rw(n851_o),
    .ctrl_i_lsu_mo_we(n852_o),
    .ctrl_i_lsu_fence(n853_o),
    .ctrl_i_lsu_priv(n854_o),
    .ctrl_i_ir_funct3(n855_o),
    .ctrl_i_ir_funct12(n856_o),
    .ctrl_i_ir_opcode(n857_o),
    .ctrl_i_cpu_priv(n858_o),
    .ctrl_i_cpu_sleep(n859_o),
    .ctrl_i_cpu_trap(n860_o),
    .ctrl_i_cpu_debug(n861_o),
    .addr_i(alu_add),
    .wdata_i(rs2),
    .pmp_fault_i(pmp_rw_fault),
    .bus_rsp_i_data(n871_o),
    .bus_rsp_i_ack(n872_o),
    .bus_rsp_i_err(n873_o),
    .rdata_o(neorv32_cpu_lsu_inst_rdata_o),
    .mar_o(neorv32_cpu_lsu_inst_mar_o),
    .wait_o(neorv32_cpu_lsu_inst_wait_o),
    .ma_load_o(neorv32_cpu_lsu_inst_ma_load_o),
    .ma_store_o(neorv32_cpu_lsu_inst_ma_store_o),
    .be_load_o(neorv32_cpu_lsu_inst_be_load_o),
    .be_store_o(neorv32_cpu_lsu_inst_be_store_o),
    .bus_req_o_addr(neorv32_cpu_lsu_inst_bus_req_o_addr),
    .bus_req_o_data(neorv32_cpu_lsu_inst_bus_req_o_data),
    .bus_req_o_ben(neorv32_cpu_lsu_inst_bus_req_o_ben),
    .bus_req_o_stb(neorv32_cpu_lsu_inst_bus_req_o_stb),
    .bus_req_o_rw(neorv32_cpu_lsu_inst_bus_req_o_rw),
    .bus_req_o_src(neorv32_cpu_lsu_inst_bus_req_o_src),
    .bus_req_o_priv(neorv32_cpu_lsu_inst_bus_req_o_priv),
    .bus_req_o_rvso(neorv32_cpu_lsu_inst_bus_req_o_rvso),
    .bus_req_o_fence(neorv32_cpu_lsu_inst_bus_req_o_fence));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:488:48  */
  assign n838_o = ctrl[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:488:62  */
  assign n839_o = ctrl[5:1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:488:38  */
  assign n840_o = ctrl[10:6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:487:43  */
  assign n841_o = ctrl[15:11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:487:48  */
  assign n842_o = ctrl[20:16]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:487:62  */
  assign n843_o = ctrl[22:21]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:487:38  */
  assign n844_o = ctrl[23]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:486:43  */
  assign n845_o = ctrl[26:24]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:486:48  */
  assign n846_o = ctrl[27]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:486:62  */
  assign n847_o = ctrl[28]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:486:38  */
  assign n848_o = ctrl[29]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:485:43  */
  assign n849_o = ctrl[35:30]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:485:48  */
  assign n850_o = ctrl[36]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:485:62  */
  assign n851_o = ctrl[37]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:485:38  */
  assign n852_o = ctrl[38]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:484:43  */
  assign n853_o = ctrl[39]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:484:48  */
  assign n854_o = ctrl[40]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:484:62  */
  assign n855_o = ctrl[43:41]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:484:38  */
  assign n856_o = ctrl[55:44]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:483:43  */
  assign n857_o = ctrl[62:56]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:483:48  */
  assign n858_o = ctrl[63]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:483:62  */
  assign n859_o = ctrl[64]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:483:38  */
  assign n860_o = ctrl[65]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:482:43  */
  assign n861_o = ctrl[66]; // extract
  assign n869_o = {neorv32_cpu_lsu_inst_bus_req_o_fence, neorv32_cpu_lsu_inst_bus_req_o_rvso, neorv32_cpu_lsu_inst_bus_req_o_priv, neorv32_cpu_lsu_inst_bus_req_o_src, neorv32_cpu_lsu_inst_bus_req_o_rw, neorv32_cpu_lsu_inst_bus_req_o_stb, neorv32_cpu_lsu_inst_bus_req_o_ben, neorv32_cpu_lsu_inst_bus_req_o_data, neorv32_cpu_lsu_inst_bus_req_o_addr};
  assign n871_o = n742_o[31:0]; // extract
  assign n872_o = n742_o[32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:471:9  */
  assign n873_o = n742_o[33]; // extract
endmodule

module neorv32_top_0_0_4_0_64_4_16384_8192_4_64_4_64_1024_32_32_8_256_0_0_1_1_1_1_1_1_0_1_32_32_1_1_1_ba529af7aa7a6f941b636046ab20a941c3aa1b01
  (input  clk_i,
   input  rstn_i,
   input  jtag_trst_i,
   input  jtag_tck_i,
   input  jtag_tdi_i,
   input  jtag_tms_i,
   input  [31:0] xbus_dat_i,
   input  xbus_ack_i,
   input  xbus_err_i,
   input  [31:0] slink_rx_dat_i,
   input  slink_rx_val_i,
   input  slink_rx_lst_i,
   input  slink_tx_rdy_i,
   input  xip_dat_i,
   input  [63:0] gpio_i,
   input  uart0_rxd_i,
   input  uart0_cts_i,
   input  uart1_rxd_i,
   input  uart1_cts_i,
   input  spi_dat_i,
   input  sdi_clk_i,
   input  sdi_dat_i,
   input  sdi_csn_i,
   input  twi_sda_i,
   input  twi_scl_i,
   input  onewire_i,
   input  [31:0] cfs_in_i,
   input  gptmr_trig_i,
   input  [31:0] xirq_i,
   input  mtime_irq_i,
   input  msw_irq_i,
   input  mext_irq_i,
   output jtag_tdo_o,
   output [31:0] xbus_adr_o,
   output [31:0] xbus_dat_o,
   output xbus_we_o,
   output [3:0] xbus_sel_o,
   output xbus_stb_o,
   output xbus_cyc_o,
   output slink_rx_rdy_o,
   output [31:0] slink_tx_dat_o,
   output slink_tx_val_o,
   output slink_tx_lst_o,
   output xip_csn_o,
   output xip_clk_o,
   output xip_dat_o,
   output [63:0] gpio_o,
   output uart0_txd_o,
   output uart0_rts_o,
   output uart1_txd_o,
   output uart1_rts_o,
   output spi_clk_o,
   output spi_dat_o,
   output [7:0] spi_csn_o,
   output sdi_dat_o,
   output twi_sda_o,
   output twi_scl_o,
   output onewire_o,
   output [11:0] pwm_o,
   output [31:0] cfs_out_o,
   output neoled_o,
   output [63:0] mtime_time_o);
  wire rstn_wdt;
  wire [3:0] rstn_sys_sreg;
  wire rstn_sys;
  wire clk_cpu;
  wire dci_ndmrstn;
  wire dci_halt_req;
  wire [73:0] cpu_i_req;
  wire [73:0] cpu_d_req;
  wire [33:0] cpu_i_rsp;
  wire [33:0] cpu_d_rsp;
  wire [73:0] icache_req;
  wire [73:0] dcache_req;
  wire [33:0] icache_rsp;
  wire [33:0] dcache_rsp;
  wire [73:0] core_req;
  wire [33:0] core_rsp;
  wire [73:0] main_req;
  wire [73:0] main2_req;
  wire [33:0] main_rsp;
  wire [33:0] main2_rsp;
  wire [73:0] io_req;
  wire [73:0] xcache_req;
  wire [73:0] xbus_req;
  wire [33:0] imem_rsp;
  wire [33:0] dmem_rsp;
  wire [33:0] xip_rsp;
  wire [33:0] boot_rsp;
  wire [33:0] io_rsp;
  wire [33:0] xcache_rsp;
  wire [33:0] xbus_rsp;
  wire [1553:0] iodev_req;
  wire [713:0] iodev_rsp;
  wire [15:0] firq;
  wire [15:0] cpu_firq;
  wire mtime_irq;
  wire [63:0] mtime_time;
  wire n197_o;
  wire n218_o;
  wire n219_o;
  wire n220_o;
  wire [2:0] n221_o;
  wire [3:0] n223_o;
  wire [3:0] n225_o;
  wire n232_o;
  wire n234_o;
  wire n236_o;
  wire n237_o;
  wire n238_o;
  wire n239_o;
  wire n240_o;
  wire n241_o;
  wire core_complex_neorv32_cpu_inst_sleep_o;
  wire core_complex_neorv32_cpu_inst_debug_o;
  wire [31:0] core_complex_neorv32_cpu_inst_ibus_req_o_addr;
  wire [31:0] core_complex_neorv32_cpu_inst_ibus_req_o_data;
  wire [3:0] core_complex_neorv32_cpu_inst_ibus_req_o_ben;
  wire core_complex_neorv32_cpu_inst_ibus_req_o_stb;
  wire core_complex_neorv32_cpu_inst_ibus_req_o_rw;
  wire core_complex_neorv32_cpu_inst_ibus_req_o_src;
  wire core_complex_neorv32_cpu_inst_ibus_req_o_priv;
  wire core_complex_neorv32_cpu_inst_ibus_req_o_rvso;
  wire core_complex_neorv32_cpu_inst_ibus_req_o_fence;
  wire [31:0] core_complex_neorv32_cpu_inst_dbus_req_o_addr;
  wire [31:0] core_complex_neorv32_cpu_inst_dbus_req_o_data;
  wire [3:0] core_complex_neorv32_cpu_inst_dbus_req_o_ben;
  wire core_complex_neorv32_cpu_inst_dbus_req_o_stb;
  wire core_complex_neorv32_cpu_inst_dbus_req_o_rw;
  wire core_complex_neorv32_cpu_inst_dbus_req_o_src;
  wire core_complex_neorv32_cpu_inst_dbus_req_o_priv;
  wire core_complex_neorv32_cpu_inst_dbus_req_o_rvso;
  wire core_complex_neorv32_cpu_inst_dbus_req_o_fence;
  wire [73:0] n340_o;
  wire [31:0] n342_o;
  wire n343_o;
  wire n344_o;
  wire [73:0] n345_o;
  wire [31:0] n347_o;
  wire n348_o;
  wire n349_o;
  wire n350_o;
  wire n351_o;
  wire n352_o;
  wire n353_o;
  wire n354_o;
  wire n355_o;
  wire n356_o;
  wire n357_o;
  wire n358_o;
  wire n359_o;
  wire n360_o;
  wire n361_o;
  wire n362_o;
  wire n363_o;
  wire n364_o;
  wire n365_o;
  wire [31:0] core_complex_neorv32_core_bus_switch_inst_a_rsp_o_data;
  wire core_complex_neorv32_core_bus_switch_inst_a_rsp_o_ack;
  wire core_complex_neorv32_core_bus_switch_inst_a_rsp_o_err;
  wire [31:0] core_complex_neorv32_core_bus_switch_inst_b_rsp_o_data;
  wire core_complex_neorv32_core_bus_switch_inst_b_rsp_o_ack;
  wire core_complex_neorv32_core_bus_switch_inst_b_rsp_o_err;
  wire [31:0] core_complex_neorv32_core_bus_switch_inst_x_req_o_addr;
  wire [31:0] core_complex_neorv32_core_bus_switch_inst_x_req_o_data;
  wire [3:0] core_complex_neorv32_core_bus_switch_inst_x_req_o_ben;
  wire core_complex_neorv32_core_bus_switch_inst_x_req_o_stb;
  wire core_complex_neorv32_core_bus_switch_inst_x_req_o_rw;
  wire core_complex_neorv32_core_bus_switch_inst_x_req_o_src;
  wire core_complex_neorv32_core_bus_switch_inst_x_req_o_priv;
  wire core_complex_neorv32_core_bus_switch_inst_x_req_o_rvso;
  wire core_complex_neorv32_core_bus_switch_inst_x_req_o_fence;
  wire [31:0] n366_o;
  wire [31:0] n367_o;
  wire [3:0] n368_o;
  wire n369_o;
  wire n370_o;
  wire n371_o;
  wire n372_o;
  wire n373_o;
  wire n374_o;
  wire [33:0] n375_o;
  wire [31:0] n377_o;
  wire [31:0] n378_o;
  wire [3:0] n379_o;
  wire n380_o;
  wire n381_o;
  wire n382_o;
  wire n383_o;
  wire n384_o;
  wire n385_o;
  wire [33:0] n386_o;
  wire [73:0] n388_o;
  wire [31:0] n390_o;
  wire n391_o;
  wire n392_o;
  wire [31:0] neorv32_bus_gateway_inst_main_rsp_o_data;
  wire neorv32_bus_gateway_inst_main_rsp_o_ack;
  wire neorv32_bus_gateway_inst_main_rsp_o_err;
  wire [31:0] neorv32_bus_gateway_inst_imem_req_o_addr;
  wire [31:0] neorv32_bus_gateway_inst_imem_req_o_data;
  wire [3:0] neorv32_bus_gateway_inst_imem_req_o_ben;
  wire neorv32_bus_gateway_inst_imem_req_o_stb;
  wire neorv32_bus_gateway_inst_imem_req_o_rw;
  wire neorv32_bus_gateway_inst_imem_req_o_src;
  wire neorv32_bus_gateway_inst_imem_req_o_priv;
  wire neorv32_bus_gateway_inst_imem_req_o_rvso;
  wire neorv32_bus_gateway_inst_imem_req_o_fence;
  wire [31:0] neorv32_bus_gateway_inst_dmem_req_o_addr;
  wire [31:0] neorv32_bus_gateway_inst_dmem_req_o_data;
  wire [3:0] neorv32_bus_gateway_inst_dmem_req_o_ben;
  wire neorv32_bus_gateway_inst_dmem_req_o_stb;
  wire neorv32_bus_gateway_inst_dmem_req_o_rw;
  wire neorv32_bus_gateway_inst_dmem_req_o_src;
  wire neorv32_bus_gateway_inst_dmem_req_o_priv;
  wire neorv32_bus_gateway_inst_dmem_req_o_rvso;
  wire neorv32_bus_gateway_inst_dmem_req_o_fence;
  wire [31:0] neorv32_bus_gateway_inst_xip_req_o_addr;
  wire [31:0] neorv32_bus_gateway_inst_xip_req_o_data;
  wire [3:0] neorv32_bus_gateway_inst_xip_req_o_ben;
  wire neorv32_bus_gateway_inst_xip_req_o_stb;
  wire neorv32_bus_gateway_inst_xip_req_o_rw;
  wire neorv32_bus_gateway_inst_xip_req_o_src;
  wire neorv32_bus_gateway_inst_xip_req_o_priv;
  wire neorv32_bus_gateway_inst_xip_req_o_rvso;
  wire neorv32_bus_gateway_inst_xip_req_o_fence;
  wire [31:0] neorv32_bus_gateway_inst_boot_req_o_addr;
  wire [31:0] neorv32_bus_gateway_inst_boot_req_o_data;
  wire [3:0] neorv32_bus_gateway_inst_boot_req_o_ben;
  wire neorv32_bus_gateway_inst_boot_req_o_stb;
  wire neorv32_bus_gateway_inst_boot_req_o_rw;
  wire neorv32_bus_gateway_inst_boot_req_o_src;
  wire neorv32_bus_gateway_inst_boot_req_o_priv;
  wire neorv32_bus_gateway_inst_boot_req_o_rvso;
  wire neorv32_bus_gateway_inst_boot_req_o_fence;
  wire [31:0] neorv32_bus_gateway_inst_io_req_o_addr;
  wire [31:0] neorv32_bus_gateway_inst_io_req_o_data;
  wire [3:0] neorv32_bus_gateway_inst_io_req_o_ben;
  wire neorv32_bus_gateway_inst_io_req_o_stb;
  wire neorv32_bus_gateway_inst_io_req_o_rw;
  wire neorv32_bus_gateway_inst_io_req_o_src;
  wire neorv32_bus_gateway_inst_io_req_o_priv;
  wire neorv32_bus_gateway_inst_io_req_o_rvso;
  wire neorv32_bus_gateway_inst_io_req_o_fence;
  wire [31:0] neorv32_bus_gateway_inst_ext_req_o_addr;
  wire [31:0] neorv32_bus_gateway_inst_ext_req_o_data;
  wire [3:0] neorv32_bus_gateway_inst_ext_req_o_ben;
  wire neorv32_bus_gateway_inst_ext_req_o_stb;
  wire neorv32_bus_gateway_inst_ext_req_o_rw;
  wire neorv32_bus_gateway_inst_ext_req_o_src;
  wire neorv32_bus_gateway_inst_ext_req_o_priv;
  wire neorv32_bus_gateway_inst_ext_req_o_rvso;
  wire neorv32_bus_gateway_inst_ext_req_o_fence;
  wire [31:0] n395_o;
  wire [31:0] n396_o;
  wire [3:0] n397_o;
  wire n398_o;
  wire n399_o;
  wire n400_o;
  wire n401_o;
  wire n402_o;
  wire n403_o;
  wire [33:0] n404_o;
  wire [31:0] n408_o;
  wire n409_o;
  wire n410_o;
  wire [31:0] n413_o;
  wire n414_o;
  wire n415_o;
  wire [31:0] n418_o;
  wire n419_o;
  wire n420_o;
  wire [31:0] n423_o;
  wire n424_o;
  wire n425_o;
  wire [73:0] n426_o;
  wire [31:0] n428_o;
  wire n429_o;
  wire n430_o;
  wire [73:0] n431_o;
  wire [31:0] n433_o;
  wire n434_o;
  wire n435_o;
  localparam n441_o = 1'b1;
  localparam n442_o = 1'b0;
  localparam n443_o = 1'b0;
  wire [31:0] memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_data;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_ack;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_err;
  wire [31:0] memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_adr_o;
  wire [31:0] memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_dat_o;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_we_o;
  wire [3:0] memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_sel_o;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_stb_o;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_cyc_o;
  wire [31:0] n444_o;
  wire [31:0] n445_o;
  wire [3:0] n446_o;
  wire n447_o;
  wire n448_o;
  wire n449_o;
  wire n450_o;
  wire n451_o;
  wire n452_o;
  wire [33:0] n453_o;
  wire [31:0] memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_data;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_ack;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_err;
  wire [31:0] memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_addr;
  wire [31:0] memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_data;
  wire [3:0] memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_ben;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_stb;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_rw;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_src;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_priv;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_rvso;
  wire memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_fence;
  wire [31:0] n461_o;
  wire [31:0] n462_o;
  wire [3:0] n463_o;
  wire n464_o;
  wire n465_o;
  wire n466_o;
  wire n467_o;
  wire n468_o;
  wire n469_o;
  wire [33:0] n470_o;
  wire [73:0] n472_o;
  wire [31:0] n474_o;
  wire n475_o;
  wire n476_o;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_main_rsp_o_data;
  wire io_system_neorv32_bus_io_switch_inst_main_rsp_o_ack;
  wire io_system_neorv32_bus_io_switch_inst_main_rsp_o_err;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_00_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_00_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_00_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_00_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_00_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_00_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_00_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_00_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_00_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_01_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_01_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_01_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_01_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_01_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_01_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_01_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_01_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_01_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_02_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_02_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_02_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_02_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_02_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_02_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_02_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_02_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_02_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_03_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_03_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_03_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_03_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_03_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_03_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_03_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_03_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_03_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_04_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_04_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_04_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_04_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_04_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_04_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_04_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_04_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_04_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_05_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_05_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_05_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_05_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_05_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_05_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_05_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_05_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_05_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_06_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_06_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_06_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_06_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_06_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_06_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_06_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_06_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_06_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_07_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_07_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_07_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_07_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_07_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_07_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_07_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_07_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_07_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_08_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_08_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_08_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_08_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_08_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_08_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_08_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_08_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_08_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_09_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_09_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_09_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_09_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_09_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_09_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_09_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_09_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_09_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_10_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_10_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_10_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_10_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_10_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_10_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_10_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_10_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_10_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_11_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_11_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_11_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_11_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_11_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_11_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_11_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_11_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_11_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_12_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_12_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_12_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_12_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_12_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_12_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_12_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_12_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_12_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_13_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_13_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_13_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_13_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_13_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_13_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_13_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_13_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_13_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_14_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_14_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_14_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_14_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_14_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_14_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_14_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_14_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_14_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_15_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_15_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_15_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_15_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_15_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_15_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_15_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_15_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_15_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_16_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_16_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_16_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_16_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_16_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_16_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_16_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_16_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_16_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_17_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_17_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_17_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_17_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_17_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_17_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_17_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_17_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_17_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_18_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_18_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_18_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_18_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_18_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_18_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_18_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_18_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_18_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_19_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_19_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_19_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_19_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_19_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_19_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_19_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_19_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_19_req_o_fence;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_20_req_o_addr;
  wire [31:0] io_system_neorv32_bus_io_switch_inst_dev_20_req_o_data;
  wire [3:0] io_system_neorv32_bus_io_switch_inst_dev_20_req_o_ben;
  wire io_system_neorv32_bus_io_switch_inst_dev_20_req_o_stb;
  wire io_system_neorv32_bus_io_switch_inst_dev_20_req_o_rw;
  wire io_system_neorv32_bus_io_switch_inst_dev_20_req_o_src;
  wire io_system_neorv32_bus_io_switch_inst_dev_20_req_o_priv;
  wire io_system_neorv32_bus_io_switch_inst_dev_20_req_o_rvso;
  wire io_system_neorv32_bus_io_switch_inst_dev_20_req_o_fence;
  wire [31:0] n477_o;
  wire [31:0] n478_o;
  wire [3:0] n479_o;
  wire n480_o;
  wire n481_o;
  wire n482_o;
  wire n483_o;
  wire n484_o;
  wire n485_o;
  wire [33:0] n486_o;
  wire [73:0] n488_o;
  wire [33:0] n490_o;
  wire [31:0] n491_o;
  wire n492_o;
  wire n493_o;
  wire [73:0] n494_o;
  wire [33:0] n496_o;
  wire [31:0] n497_o;
  wire n498_o;
  wire n499_o;
  wire [73:0] n500_o;
  wire [33:0] n502_o;
  wire [31:0] n503_o;
  wire n504_o;
  wire n505_o;
  wire [73:0] n506_o;
  wire [33:0] n508_o;
  wire [31:0] n509_o;
  wire n510_o;
  wire n511_o;
  wire [73:0] n512_o;
  wire [33:0] n514_o;
  wire [31:0] n515_o;
  wire n516_o;
  wire n517_o;
  wire [73:0] n518_o;
  wire [33:0] n520_o;
  wire [31:0] n521_o;
  wire n522_o;
  wire n523_o;
  wire [73:0] n524_o;
  wire [33:0] n526_o;
  wire [31:0] n527_o;
  wire n528_o;
  wire n529_o;
  wire [73:0] n530_o;
  wire [33:0] n532_o;
  wire [31:0] n533_o;
  wire n534_o;
  wire n535_o;
  wire [73:0] n536_o;
  wire [33:0] n538_o;
  wire [31:0] n539_o;
  wire n540_o;
  wire n541_o;
  wire [73:0] n542_o;
  wire [33:0] n544_o;
  wire [31:0] n545_o;
  wire n546_o;
  wire n547_o;
  wire [73:0] n548_o;
  wire [33:0] n550_o;
  wire [31:0] n551_o;
  wire n552_o;
  wire n553_o;
  wire [73:0] n554_o;
  wire [33:0] n556_o;
  wire [31:0] n557_o;
  wire n558_o;
  wire n559_o;
  wire [73:0] n560_o;
  wire [33:0] n562_o;
  wire [31:0] n563_o;
  wire n564_o;
  wire n565_o;
  wire [73:0] n566_o;
  wire [33:0] n568_o;
  wire [31:0] n569_o;
  wire n570_o;
  wire n571_o;
  wire [73:0] n572_o;
  wire [33:0] n574_o;
  wire [31:0] n575_o;
  wire n576_o;
  wire n577_o;
  wire [73:0] n578_o;
  wire [33:0] n580_o;
  wire [31:0] n581_o;
  wire n582_o;
  wire n583_o;
  wire [73:0] n584_o;
  wire [33:0] n586_o;
  wire [31:0] n587_o;
  wire n588_o;
  wire n589_o;
  wire [73:0] n590_o;
  wire [33:0] n592_o;
  wire [31:0] n593_o;
  wire n594_o;
  wire n595_o;
  wire [73:0] n596_o;
  wire [33:0] n598_o;
  wire [31:0] n599_o;
  wire n600_o;
  wire n601_o;
  wire [73:0] n602_o;
  wire [33:0] n604_o;
  wire [31:0] n605_o;
  wire n606_o;
  wire n607_o;
  wire [73:0] n608_o;
  wire [33:0] n610_o;
  wire [31:0] n611_o;
  wire n612_o;
  wire n613_o;
  localparam [31:0] n616_o = 32'b00000000000000000000000000000000;
  localparam n617_o = 1'b0;
  localparam [63:0] n619_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_data;
  wire io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_ack;
  wire io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_err;
  wire [63:0] io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_time_o;
  wire io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_irq_o;
  wire [73:0] n623_o;
  wire [31:0] n624_o;
  wire [31:0] n625_o;
  wire [3:0] n626_o;
  wire n627_o;
  wire n628_o;
  wire n629_o;
  wire n630_o;
  wire n631_o;
  wire n632_o;
  wire [33:0] n633_o;
  wire n638_o;
  wire [31:0] n641_o;
  wire [31:0] n646_o;
  localparam n647_o = 1'b0;
  localparam n648_o = 1'b1;
  localparam n652_o = 1'b0;
  localparam n653_o = 1'b1;
  localparam n657_o = 1'b0;
  localparam n658_o = 1'b0;
  localparam [7:0] n659_o = 8'b11111111;
  localparam n662_o = 1'b1;
  localparam n663_o = 1'b1;
  localparam [11:0] n667_o = 12'b000000000000;
  localparam n671_o = 1'b0;
  localparam n675_o = 1'b1;
  localparam n679_o = 1'b0;
  localparam [31:0] n680_o = 32'b00000000000000000000000000000000;
  localparam n681_o = 1'b0;
  localparam n682_o = 1'b0;
  wire [31:0] io_system_neorv32_sysinfo_inst_bus_rsp_o_data;
  wire io_system_neorv32_sysinfo_inst_bus_rsp_o_ack;
  wire io_system_neorv32_sysinfo_inst_bus_rsp_o_err;
  wire [73:0] n683_o;
  wire [31:0] n684_o;
  wire [31:0] n685_o;
  wire [3:0] n686_o;
  wire n687_o;
  wire n688_o;
  wire n689_o;
  wire n690_o;
  wire n691_o;
  wire n692_o;
  wire [33:0] n693_o;
  reg [3:0] n697_q;
  reg n699_q;
  wire [1553:0] n713_o;
  wire [713:0] n714_o;
  wire [15:0] n715_o;
  wire [15:0] n716_o;
  reg [31:0] n717_q;
  wire [63:0] n718_o;
  assign jtag_tdo_o = jtag_tdi_i; //(module output)
  assign xbus_adr_o = memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_adr_o; //(module output)
  assign xbus_dat_o = memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_dat_o; //(module output)
  assign xbus_we_o = memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_we_o; //(module output)
  assign xbus_sel_o = memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_sel_o; //(module output)
  assign xbus_stb_o = memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_stb_o; //(module output)
  assign xbus_cyc_o = memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_cyc_o; //(module output)
  assign slink_rx_rdy_o = n679_o; //(module output)
  assign slink_tx_dat_o = n680_o; //(module output)
  assign slink_tx_val_o = n681_o; //(module output)
  assign slink_tx_lst_o = n682_o; //(module output)
  assign xip_csn_o = n441_o; //(module output)
  assign xip_clk_o = n442_o; //(module output)
  assign xip_dat_o = n443_o; //(module output)
  assign gpio_o = n619_o; //(module output)
  assign uart0_txd_o = n647_o; //(module output)
  assign uart0_rts_o = n648_o; //(module output)
  assign uart1_txd_o = n652_o; //(module output)
  assign uart1_rts_o = n653_o; //(module output)
  assign spi_clk_o = n657_o; //(module output)
  assign spi_dat_o = n658_o; //(module output)
  assign spi_csn_o = n659_o; //(module output)
  assign sdi_dat_o = n617_o; //(module output)
  assign twi_sda_o = n662_o; //(module output)
  assign twi_scl_o = n663_o; //(module output)
  assign onewire_o = n675_o; //(module output)
  assign pwm_o = n667_o; //(module output)
  assign cfs_out_o = n616_o; //(module output)
  assign neoled_o = n671_o; //(module output)
  assign mtime_time_o = n718_o; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:288:10  */
  assign rstn_wdt = 1'b1; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:289:10  */
  assign rstn_sys_sreg = n697_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:290:10  */
  assign rstn_sys = n699_q; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:294:10  */
  assign clk_cpu = clk_i; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:313:10  */
  assign dci_ndmrstn = 1'b1; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:313:23  */
  assign dci_halt_req = 1'b0; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:316:10  */
  assign cpu_i_req = n340_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:316:22  */
  assign cpu_d_req = n345_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:317:10  */
  assign cpu_i_rsp = icache_rsp; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:317:22  */
  assign cpu_d_rsp = dcache_rsp; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:318:10  */
  assign icache_req = cpu_i_req; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:318:22  */
  assign dcache_req = cpu_d_req; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:319:10  */
  assign icache_rsp = n386_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:319:22  */
  assign dcache_rsp = n375_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:320:10  */
  assign core_req = n388_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:321:10  */
  assign core_rsp = main_rsp; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:324:10  */
  assign main_req = core_req; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:324:20  */
  assign main2_req = main_req; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:325:10  */
  assign main_rsp = main2_rsp; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:325:20  */
  assign main2_rsp = n404_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:328:63  */
  assign io_req = n426_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:328:71  */
  assign xcache_req = n472_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:328:83  */
  assign xbus_req = n431_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:329:10  */
  assign imem_rsp = 34'b0000000000000000000000000000000000; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:329:20  */
  assign dmem_rsp = 34'b0000000000000000000000000000000000; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:329:44  */
  assign xip_rsp = 34'b0000000000000000000000000000000000; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:329:53  */
  assign boot_rsp = 34'b0000000000000000000000000000000000; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:329:63  */
  assign io_rsp = n486_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:329:71  */
  assign xcache_rsp = n453_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:329:83  */
  assign xbus_rsp = n470_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:339:10  */
  assign iodev_req = n713_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:340:10  */
  assign iodev_rsp = n714_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:348:10  */
  assign firq = n715_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:349:10  */
  assign cpu_firq = n716_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:350:10  */
  assign mtime_irq = io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_irq_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:353:10  */
  assign mtime_time = io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_time_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:425:18  */
  assign n197_o = ~rstn_i;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:435:22  */
  assign n218_o = ~rstn_wdt;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:435:45  */
  assign n219_o = ~dci_ndmrstn;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:435:29  */
  assign n220_o = n218_o | n219_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:438:41  */
  assign n221_o = rstn_sys_sreg[2:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:438:73  */
  assign n223_o = {n221_o, 1'b1};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:435:9  */
  assign n225_o = n220_o ? 4'b0000 : n223_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n232_o = rstn_sys_sreg[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n234_o = 1'b1 & n232_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n236_o = rstn_sys_sreg[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n237_o = n234_o & n236_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n238_o = rstn_sys_sreg[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n239_o = n237_o & n238_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:31  */
  assign n240_o = rstn_sys_sreg[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_package.vhd:1038:22  */
  assign n241_o = n239_o & n240_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:525:5  */
  neorv32_cpu_0_4_0_64_16973a3472ca3522cdc18159c73abb10ac4c9817 core_complex_neorv32_cpu_inst (
    .clk_i(clk_cpu),
    .clk_aux_i(clk_i),
    .rstn_i(rstn_sys),
    .msi_i(msw_irq_i),
    .mei_i(mext_irq_i),
    .mti_i(mtime_irq),
    .firq_i(cpu_firq),
    .dbi_i(dci_halt_req),
    .ibus_rsp_i_data(n342_o),
    .ibus_rsp_i_ack(n343_o),
    .ibus_rsp_i_err(n344_o),
    .dbus_rsp_i_data(n347_o),
    .dbus_rsp_i_ack(n348_o),
    .dbus_rsp_i_err(n349_o),
    .sleep_o(),
    .debug_o(),
    .ibus_req_o_addr(core_complex_neorv32_cpu_inst_ibus_req_o_addr),
    .ibus_req_o_data(core_complex_neorv32_cpu_inst_ibus_req_o_data),
    .ibus_req_o_ben(core_complex_neorv32_cpu_inst_ibus_req_o_ben),
    .ibus_req_o_stb(core_complex_neorv32_cpu_inst_ibus_req_o_stb),
    .ibus_req_o_rw(core_complex_neorv32_cpu_inst_ibus_req_o_rw),
    .ibus_req_o_src(core_complex_neorv32_cpu_inst_ibus_req_o_src),
    .ibus_req_o_priv(core_complex_neorv32_cpu_inst_ibus_req_o_priv),
    .ibus_req_o_rvso(core_complex_neorv32_cpu_inst_ibus_req_o_rvso),
    .ibus_req_o_fence(core_complex_neorv32_cpu_inst_ibus_req_o_fence),
    .dbus_req_o_addr(core_complex_neorv32_cpu_inst_dbus_req_o_addr),
    .dbus_req_o_data(core_complex_neorv32_cpu_inst_dbus_req_o_data),
    .dbus_req_o_ben(core_complex_neorv32_cpu_inst_dbus_req_o_ben),
    .dbus_req_o_stb(core_complex_neorv32_cpu_inst_dbus_req_o_stb),
    .dbus_req_o_rw(core_complex_neorv32_cpu_inst_dbus_req_o_rw),
    .dbus_req_o_src(core_complex_neorv32_cpu_inst_dbus_req_o_src),
    .dbus_req_o_priv(core_complex_neorv32_cpu_inst_dbus_req_o_priv),
    .dbus_req_o_rvso(core_complex_neorv32_cpu_inst_dbus_req_o_rvso),
    .dbus_req_o_fence(core_complex_neorv32_cpu_inst_dbus_req_o_fence));
  assign n340_o = {core_complex_neorv32_cpu_inst_ibus_req_o_fence, core_complex_neorv32_cpu_inst_ibus_req_o_rvso, core_complex_neorv32_cpu_inst_ibus_req_o_priv, core_complex_neorv32_cpu_inst_ibus_req_o_src, core_complex_neorv32_cpu_inst_ibus_req_o_rw, core_complex_neorv32_cpu_inst_ibus_req_o_stb, core_complex_neorv32_cpu_inst_ibus_req_o_ben, core_complex_neorv32_cpu_inst_ibus_req_o_data, core_complex_neorv32_cpu_inst_ibus_req_o_addr};
  assign n342_o = cpu_i_rsp[31:0]; // extract
  assign n343_o = cpu_i_rsp[32]; // extract
  assign n344_o = cpu_i_rsp[33]; // extract
  assign n345_o = {core_complex_neorv32_cpu_inst_dbus_req_o_fence, core_complex_neorv32_cpu_inst_dbus_req_o_rvso, core_complex_neorv32_cpu_inst_dbus_req_o_priv, core_complex_neorv32_cpu_inst_dbus_req_o_src, core_complex_neorv32_cpu_inst_dbus_req_o_rw, core_complex_neorv32_cpu_inst_dbus_req_o_stb, core_complex_neorv32_cpu_inst_dbus_req_o_ben, core_complex_neorv32_cpu_inst_dbus_req_o_data, core_complex_neorv32_cpu_inst_dbus_req_o_addr};
  assign n347_o = cpu_d_rsp[31:0]; // extract
  assign n348_o = cpu_d_rsp[32]; // extract
  assign n349_o = cpu_d_rsp[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:584:25  */
  assign n350_o = firq[15]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:585:25  */
  assign n351_o = firq[7]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:586:25  */
  assign n352_o = firq[14]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:587:25  */
  assign n353_o = firq[13]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:588:25  */
  assign n354_o = firq[12]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:589:25  */
  assign n355_o = firq[11]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:590:25  */
  assign n356_o = firq[10]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:591:25  */
  assign n357_o = firq[8]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:592:25  */
  assign n358_o = firq[5]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:593:25  */
  assign n359_o = firq[6]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:594:25  */
  assign n360_o = firq[2]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:595:25  */
  assign n361_o = firq[9]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:596:25  */
  assign n362_o = firq[4]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:597:25  */
  assign n363_o = firq[3]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:598:25  */
  assign n364_o = firq[0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:599:25  */
  assign n365_o = firq[1]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:662:5  */
  neorv32_bus_switch_3f29546453678b855931c174a97d6c0894b8f546 core_complex_neorv32_core_bus_switch_inst (
    .clk_i(clk_cpu),
    .rstn_i(rstn_sys),
    .a_req_i_addr(n366_o),
    .a_req_i_data(n367_o),
    .a_req_i_ben(n368_o),
    .a_req_i_stb(n369_o),
    .a_req_i_rw(n370_o),
    .a_req_i_src(n371_o),
    .a_req_i_priv(n372_o),
    .a_req_i_rvso(n373_o),
    .a_req_i_fence(n374_o),
    .b_req_i_addr(n377_o),
    .b_req_i_data(n378_o),
    .b_req_i_ben(n379_o),
    .b_req_i_stb(n380_o),
    .b_req_i_rw(n381_o),
    .b_req_i_src(n382_o),
    .b_req_i_priv(n383_o),
    .b_req_i_rvso(n384_o),
    .b_req_i_fence(n385_o),
    .x_rsp_i_data(n390_o),
    .x_rsp_i_ack(n391_o),
    .x_rsp_i_err(n392_o),
    .a_rsp_o_data(core_complex_neorv32_core_bus_switch_inst_a_rsp_o_data),
    .a_rsp_o_ack(core_complex_neorv32_core_bus_switch_inst_a_rsp_o_ack),
    .a_rsp_o_err(core_complex_neorv32_core_bus_switch_inst_a_rsp_o_err),
    .b_rsp_o_data(core_complex_neorv32_core_bus_switch_inst_b_rsp_o_data),
    .b_rsp_o_ack(core_complex_neorv32_core_bus_switch_inst_b_rsp_o_ack),
    .b_rsp_o_err(core_complex_neorv32_core_bus_switch_inst_b_rsp_o_err),
    .x_req_o_addr(core_complex_neorv32_core_bus_switch_inst_x_req_o_addr),
    .x_req_o_data(core_complex_neorv32_core_bus_switch_inst_x_req_o_data),
    .x_req_o_ben(core_complex_neorv32_core_bus_switch_inst_x_req_o_ben),
    .x_req_o_stb(core_complex_neorv32_core_bus_switch_inst_x_req_o_stb),
    .x_req_o_rw(core_complex_neorv32_core_bus_switch_inst_x_req_o_rw),
    .x_req_o_src(core_complex_neorv32_core_bus_switch_inst_x_req_o_src),
    .x_req_o_priv(core_complex_neorv32_core_bus_switch_inst_x_req_o_priv),
    .x_req_o_rvso(core_complex_neorv32_core_bus_switch_inst_x_req_o_rvso),
    .x_req_o_fence(core_complex_neorv32_core_bus_switch_inst_x_req_o_fence));
  assign n366_o = dcache_req[31:0]; // extract
  assign n367_o = dcache_req[63:32]; // extract
  assign n368_o = dcache_req[67:64]; // extract
  assign n369_o = dcache_req[68]; // extract
  assign n370_o = dcache_req[69]; // extract
  assign n371_o = dcache_req[70]; // extract
  assign n372_o = dcache_req[71]; // extract
  assign n373_o = dcache_req[72]; // extract
  assign n374_o = dcache_req[73]; // extract
  assign n375_o = {core_complex_neorv32_core_bus_switch_inst_a_rsp_o_err, core_complex_neorv32_core_bus_switch_inst_a_rsp_o_ack, core_complex_neorv32_core_bus_switch_inst_a_rsp_o_data};
  assign n377_o = icache_req[31:0]; // extract
  assign n378_o = icache_req[63:32]; // extract
  assign n379_o = icache_req[67:64]; // extract
  assign n380_o = icache_req[68]; // extract
  assign n381_o = icache_req[69]; // extract
  assign n382_o = icache_req[70]; // extract
  assign n383_o = icache_req[71]; // extract
  assign n384_o = icache_req[72]; // extract
  assign n385_o = icache_req[73]; // extract
  assign n386_o = {core_complex_neorv32_core_bus_switch_inst_b_rsp_o_err, core_complex_neorv32_core_bus_switch_inst_b_rsp_o_ack, core_complex_neorv32_core_bus_switch_inst_b_rsp_o_data};
  assign n388_o = {core_complex_neorv32_core_bus_switch_inst_x_req_o_fence, core_complex_neorv32_core_bus_switch_inst_x_req_o_rvso, core_complex_neorv32_core_bus_switch_inst_x_req_o_priv, core_complex_neorv32_core_bus_switch_inst_x_req_o_src, core_complex_neorv32_core_bus_switch_inst_x_req_o_rw, core_complex_neorv32_core_bus_switch_inst_x_req_o_stb, core_complex_neorv32_core_bus_switch_inst_x_req_o_ben, core_complex_neorv32_core_bus_switch_inst_x_req_o_data, core_complex_neorv32_core_bus_switch_inst_x_req_o_addr};
  assign n390_o = core_rsp[31:0]; // extract
  assign n391_o = core_rsp[32]; // extract
  assign n392_o = core_rsp[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:763:3  */
  neorv32_bus_gateway_15_16384_8192_268435456_8192_8192_a510945699945b5d171ba29323e989d87bc97675 neorv32_bus_gateway_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .main_req_i_addr(n395_o),
    .main_req_i_data(n396_o),
    .main_req_i_ben(n397_o),
    .main_req_i_stb(n398_o),
    .main_req_i_rw(n399_o),
    .main_req_i_src(n400_o),
    .main_req_i_priv(n401_o),
    .main_req_i_rvso(n402_o),
    .main_req_i_fence(n403_o),
    .imem_rsp_i_data(n408_o),
    .imem_rsp_i_ack(n409_o),
    .imem_rsp_i_err(n410_o),
    .dmem_rsp_i_data(n413_o),
    .dmem_rsp_i_ack(n414_o),
    .dmem_rsp_i_err(n415_o),
    .xip_rsp_i_data(n418_o),
    .xip_rsp_i_ack(n419_o),
    .xip_rsp_i_err(n420_o),
    .boot_rsp_i_data(n423_o),
    .boot_rsp_i_ack(n424_o),
    .boot_rsp_i_err(n425_o),
    .io_rsp_i_data(n428_o),
    .io_rsp_i_ack(n429_o),
    .io_rsp_i_err(n430_o),
    .ext_rsp_i_data(n433_o),
    .ext_rsp_i_ack(n434_o),
    .ext_rsp_i_err(n435_o),
    .main_rsp_o_data(neorv32_bus_gateway_inst_main_rsp_o_data),
    .main_rsp_o_ack(neorv32_bus_gateway_inst_main_rsp_o_ack),
    .main_rsp_o_err(neorv32_bus_gateway_inst_main_rsp_o_err),
    .imem_req_o_addr(),
    .imem_req_o_data(),
    .imem_req_o_ben(),
    .imem_req_o_stb(),
    .imem_req_o_rw(),
    .imem_req_o_src(),
    .imem_req_o_priv(),
    .imem_req_o_rvso(),
    .imem_req_o_fence(),
    .dmem_req_o_addr(),
    .dmem_req_o_data(),
    .dmem_req_o_ben(),
    .dmem_req_o_stb(),
    .dmem_req_o_rw(),
    .dmem_req_o_src(),
    .dmem_req_o_priv(),
    .dmem_req_o_rvso(),
    .dmem_req_o_fence(),
    .xip_req_o_addr(),
    .xip_req_o_data(),
    .xip_req_o_ben(),
    .xip_req_o_stb(),
    .xip_req_o_rw(),
    .xip_req_o_src(),
    .xip_req_o_priv(),
    .xip_req_o_rvso(),
    .xip_req_o_fence(),
    .boot_req_o_addr(),
    .boot_req_o_data(),
    .boot_req_o_ben(),
    .boot_req_o_stb(),
    .boot_req_o_rw(),
    .boot_req_o_src(),
    .boot_req_o_priv(),
    .boot_req_o_rvso(),
    .boot_req_o_fence(),
    .io_req_o_addr(neorv32_bus_gateway_inst_io_req_o_addr),
    .io_req_o_data(neorv32_bus_gateway_inst_io_req_o_data),
    .io_req_o_ben(neorv32_bus_gateway_inst_io_req_o_ben),
    .io_req_o_stb(neorv32_bus_gateway_inst_io_req_o_stb),
    .io_req_o_rw(neorv32_bus_gateway_inst_io_req_o_rw),
    .io_req_o_src(neorv32_bus_gateway_inst_io_req_o_src),
    .io_req_o_priv(neorv32_bus_gateway_inst_io_req_o_priv),
    .io_req_o_rvso(neorv32_bus_gateway_inst_io_req_o_rvso),
    .io_req_o_fence(neorv32_bus_gateway_inst_io_req_o_fence),
    .ext_req_o_addr(neorv32_bus_gateway_inst_ext_req_o_addr),
    .ext_req_o_data(neorv32_bus_gateway_inst_ext_req_o_data),
    .ext_req_o_ben(neorv32_bus_gateway_inst_ext_req_o_ben),
    .ext_req_o_stb(neorv32_bus_gateway_inst_ext_req_o_stb),
    .ext_req_o_rw(neorv32_bus_gateway_inst_ext_req_o_rw),
    .ext_req_o_src(neorv32_bus_gateway_inst_ext_req_o_src),
    .ext_req_o_priv(neorv32_bus_gateway_inst_ext_req_o_priv),
    .ext_req_o_rvso(neorv32_bus_gateway_inst_ext_req_o_rvso),
    .ext_req_o_fence(neorv32_bus_gateway_inst_ext_req_o_fence));
  assign n395_o = main2_req[31:0]; // extract
  assign n396_o = main2_req[63:32]; // extract
  assign n397_o = main2_req[67:64]; // extract
  assign n398_o = main2_req[68]; // extract
  assign n399_o = main2_req[69]; // extract
  assign n400_o = main2_req[70]; // extract
  assign n401_o = main2_req[71]; // extract
  assign n402_o = main2_req[72]; // extract
  assign n403_o = main2_req[73]; // extract
  assign n404_o = {neorv32_bus_gateway_inst_main_rsp_o_err, neorv32_bus_gateway_inst_main_rsp_o_ack, neorv32_bus_gateway_inst_main_rsp_o_data};
  assign n408_o = imem_rsp[31:0]; // extract
  assign n409_o = imem_rsp[32]; // extract
  assign n410_o = imem_rsp[33]; // extract
  assign n413_o = dmem_rsp[31:0]; // extract
  assign n414_o = dmem_rsp[32]; // extract
  assign n415_o = dmem_rsp[33]; // extract
  assign n418_o = xip_rsp[31:0]; // extract
  assign n419_o = xip_rsp[32]; // extract
  assign n420_o = xip_rsp[33]; // extract
  assign n423_o = boot_rsp[31:0]; // extract
  assign n424_o = boot_rsp[32]; // extract
  assign n425_o = boot_rsp[33]; // extract
  assign n426_o = {neorv32_bus_gateway_inst_io_req_o_fence, neorv32_bus_gateway_inst_io_req_o_rvso, neorv32_bus_gateway_inst_io_req_o_priv, neorv32_bus_gateway_inst_io_req_o_src, neorv32_bus_gateway_inst_io_req_o_rw, neorv32_bus_gateway_inst_io_req_o_stb, neorv32_bus_gateway_inst_io_req_o_ben, neorv32_bus_gateway_inst_io_req_o_data, neorv32_bus_gateway_inst_io_req_o_addr};
  assign n428_o = io_rsp[31:0]; // extract
  assign n429_o = io_rsp[32]; // extract
  assign n430_o = io_rsp[33]; // extract
  assign n431_o = {neorv32_bus_gateway_inst_ext_req_o_fence, neorv32_bus_gateway_inst_ext_req_o_rvso, neorv32_bus_gateway_inst_ext_req_o_priv, neorv32_bus_gateway_inst_ext_req_o_src, neorv32_bus_gateway_inst_ext_req_o_rw, neorv32_bus_gateway_inst_ext_req_o_stb, neorv32_bus_gateway_inst_ext_req_o_ben, neorv32_bus_gateway_inst_ext_req_o_data, neorv32_bus_gateway_inst_ext_req_o_addr};
  assign n433_o = xbus_rsp[31:0]; // extract
  assign n434_o = xbus_rsp[32]; // extract
  assign n435_o = xbus_rsp[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:953:7  */
  neorv32_xbus_1024_eee447edc79fea1ca7c7d34e463261cda4ba339e memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .bus_req_i_addr(n444_o),
    .bus_req_i_data(n445_o),
    .bus_req_i_ben(n446_o),
    .bus_req_i_stb(n447_o),
    .bus_req_i_rw(n448_o),
    .bus_req_i_src(n449_o),
    .bus_req_i_priv(n450_o),
    .bus_req_i_rvso(n451_o),
    .bus_req_i_fence(n452_o),
    .xbus_dat_i(xbus_dat_i),
    .xbus_ack_i(xbus_ack_i),
    .xbus_err_i(xbus_err_i),
    .bus_rsp_o_data(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_data),
    .bus_rsp_o_ack(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_ack),
    .bus_rsp_o_err(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_err),
    .xbus_adr_o(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_adr_o),
    .xbus_dat_o(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_dat_o),
    .xbus_we_o(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_we_o),
    .xbus_sel_o(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_sel_o),
    .xbus_stb_o(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_stb_o),
    .xbus_cyc_o(memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_xbus_cyc_o));
  assign n444_o = xcache_req[31:0]; // extract
  assign n445_o = xcache_req[63:32]; // extract
  assign n446_o = xcache_req[67:64]; // extract
  assign n447_o = xcache_req[68]; // extract
  assign n448_o = xcache_req[69]; // extract
  assign n449_o = xcache_req[70]; // extract
  assign n450_o = xcache_req[71]; // extract
  assign n451_o = xcache_req[72]; // extract
  assign n452_o = xcache_req[73]; // extract
  assign n453_o = {memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_err, memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_ack, memory_system_neorv32_xbus_inst_true_neorv32_xbus_inst_bus_rsp_o_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:980:9  */
  neorv32_cache_32_32_b2a9daee4605f0af85049a2738d2ab5c0686fc65 memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .host_req_i_addr(n461_o),
    .host_req_i_data(n462_o),
    .host_req_i_ben(n463_o),
    .host_req_i_stb(n464_o),
    .host_req_i_rw(n465_o),
    .host_req_i_src(n466_o),
    .host_req_i_priv(n467_o),
    .host_req_i_rvso(n468_o),
    .host_req_i_fence(n469_o),
    .bus_rsp_i_data(n474_o),
    .bus_rsp_i_ack(n475_o),
    .bus_rsp_i_err(n476_o),
    .host_rsp_o_data(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_data),
    .host_rsp_o_ack(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_ack),
    .host_rsp_o_err(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_err),
    .bus_req_o_addr(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_addr),
    .bus_req_o_data(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_data),
    .bus_req_o_ben(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_ben),
    .bus_req_o_stb(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_stb),
    .bus_req_o_rw(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_rw),
    .bus_req_o_src(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_src),
    .bus_req_o_priv(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_priv),
    .bus_req_o_rvso(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_rvso),
    .bus_req_o_fence(memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_fence));
  assign n461_o = xbus_req[31:0]; // extract
  assign n462_o = xbus_req[63:32]; // extract
  assign n463_o = xbus_req[67:64]; // extract
  assign n464_o = xbus_req[68]; // extract
  assign n465_o = xbus_req[69]; // extract
  assign n466_o = xbus_req[70]; // extract
  assign n467_o = xbus_req[71]; // extract
  assign n468_o = xbus_req[72]; // extract
  assign n469_o = xbus_req[73]; // extract
  assign n470_o = {memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_err, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_ack, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_host_rsp_o_data};
  assign n472_o = {memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_fence, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_rvso, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_priv, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_src, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_rw, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_stb, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_ben, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_data, memory_system_neorv32_xbus_inst_true_neorv32_xcache_inst_true_neorv32_xcache_inst_bus_req_o_addr};
  assign n474_o = xcache_rsp[31:0]; // extract
  assign n475_o = xcache_rsp[32]; // extract
  assign n476_o = xcache_rsp[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1028:5  */
  neorv32_bus_io_switch_256_84bc3e102e5c7d00d4cf85e98418cab7f8480bb6 io_system_neorv32_bus_io_switch_inst (
    .main_req_i_addr(n477_o),
    .main_req_i_data(n478_o),
    .main_req_i_ben(n479_o),
    .main_req_i_stb(n480_o),
    .main_req_i_rw(n481_o),
    .main_req_i_src(n482_o),
    .main_req_i_priv(n483_o),
    .main_req_i_rvso(n484_o),
    .main_req_i_fence(n485_o),
    .dev_00_rsp_i_data(n491_o),
    .dev_00_rsp_i_ack(n492_o),
    .dev_00_rsp_i_err(n493_o),
    .dev_01_rsp_i_data(n497_o),
    .dev_01_rsp_i_ack(n498_o),
    .dev_01_rsp_i_err(n499_o),
    .dev_02_rsp_i_data(n503_o),
    .dev_02_rsp_i_ack(n504_o),
    .dev_02_rsp_i_err(n505_o),
    .dev_03_rsp_i_data(n509_o),
    .dev_03_rsp_i_ack(n510_o),
    .dev_03_rsp_i_err(n511_o),
    .dev_04_rsp_i_data(n515_o),
    .dev_04_rsp_i_ack(n516_o),
    .dev_04_rsp_i_err(n517_o),
    .dev_05_rsp_i_data(n521_o),
    .dev_05_rsp_i_ack(n522_o),
    .dev_05_rsp_i_err(n523_o),
    .dev_06_rsp_i_data(n527_o),
    .dev_06_rsp_i_ack(n528_o),
    .dev_06_rsp_i_err(n529_o),
    .dev_07_rsp_i_data(n533_o),
    .dev_07_rsp_i_ack(n534_o),
    .dev_07_rsp_i_err(n535_o),
    .dev_08_rsp_i_data(n539_o),
    .dev_08_rsp_i_ack(n540_o),
    .dev_08_rsp_i_err(n541_o),
    .dev_09_rsp_i_data(n545_o),
    .dev_09_rsp_i_ack(n546_o),
    .dev_09_rsp_i_err(n547_o),
    .dev_10_rsp_i_data(n551_o),
    .dev_10_rsp_i_ack(n552_o),
    .dev_10_rsp_i_err(n553_o),
    .dev_11_rsp_i_data(n557_o),
    .dev_11_rsp_i_ack(n558_o),
    .dev_11_rsp_i_err(n559_o),
    .dev_12_rsp_i_data(n563_o),
    .dev_12_rsp_i_ack(n564_o),
    .dev_12_rsp_i_err(n565_o),
    .dev_13_rsp_i_data(n569_o),
    .dev_13_rsp_i_ack(n570_o),
    .dev_13_rsp_i_err(n571_o),
    .dev_14_rsp_i_data(n575_o),
    .dev_14_rsp_i_ack(n576_o),
    .dev_14_rsp_i_err(n577_o),
    .dev_15_rsp_i_data(n581_o),
    .dev_15_rsp_i_ack(n582_o),
    .dev_15_rsp_i_err(n583_o),
    .dev_16_rsp_i_data(n587_o),
    .dev_16_rsp_i_ack(n588_o),
    .dev_16_rsp_i_err(n589_o),
    .dev_17_rsp_i_data(n593_o),
    .dev_17_rsp_i_ack(n594_o),
    .dev_17_rsp_i_err(n595_o),
    .dev_18_rsp_i_data(n599_o),
    .dev_18_rsp_i_ack(n600_o),
    .dev_18_rsp_i_err(n601_o),
    .dev_19_rsp_i_data(n605_o),
    .dev_19_rsp_i_ack(n606_o),
    .dev_19_rsp_i_err(n607_o),
    .dev_20_rsp_i_data(n611_o),
    .dev_20_rsp_i_ack(n612_o),
    .dev_20_rsp_i_err(n613_o),
    .main_rsp_o_data(io_system_neorv32_bus_io_switch_inst_main_rsp_o_data),
    .main_rsp_o_ack(io_system_neorv32_bus_io_switch_inst_main_rsp_o_ack),
    .main_rsp_o_err(io_system_neorv32_bus_io_switch_inst_main_rsp_o_err),
    .dev_00_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_addr),
    .dev_00_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_data),
    .dev_00_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_ben),
    .dev_00_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_stb),
    .dev_00_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_rw),
    .dev_00_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_src),
    .dev_00_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_priv),
    .dev_00_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_rvso),
    .dev_00_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_00_req_o_fence),
    .dev_01_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_addr),
    .dev_01_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_data),
    .dev_01_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_ben),
    .dev_01_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_stb),
    .dev_01_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_rw),
    .dev_01_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_src),
    .dev_01_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_priv),
    .dev_01_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_rvso),
    .dev_01_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_01_req_o_fence),
    .dev_02_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_addr),
    .dev_02_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_data),
    .dev_02_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_ben),
    .dev_02_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_stb),
    .dev_02_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_rw),
    .dev_02_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_src),
    .dev_02_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_priv),
    .dev_02_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_rvso),
    .dev_02_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_02_req_o_fence),
    .dev_03_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_addr),
    .dev_03_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_data),
    .dev_03_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_ben),
    .dev_03_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_stb),
    .dev_03_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_rw),
    .dev_03_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_src),
    .dev_03_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_priv),
    .dev_03_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_rvso),
    .dev_03_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_03_req_o_fence),
    .dev_04_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_addr),
    .dev_04_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_data),
    .dev_04_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_ben),
    .dev_04_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_stb),
    .dev_04_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_rw),
    .dev_04_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_src),
    .dev_04_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_priv),
    .dev_04_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_rvso),
    .dev_04_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_04_req_o_fence),
    .dev_05_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_addr),
    .dev_05_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_data),
    .dev_05_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_ben),
    .dev_05_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_stb),
    .dev_05_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_rw),
    .dev_05_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_src),
    .dev_05_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_priv),
    .dev_05_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_rvso),
    .dev_05_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_05_req_o_fence),
    .dev_06_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_addr),
    .dev_06_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_data),
    .dev_06_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_ben),
    .dev_06_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_stb),
    .dev_06_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_rw),
    .dev_06_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_src),
    .dev_06_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_priv),
    .dev_06_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_rvso),
    .dev_06_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_06_req_o_fence),
    .dev_07_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_addr),
    .dev_07_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_data),
    .dev_07_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_ben),
    .dev_07_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_stb),
    .dev_07_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_rw),
    .dev_07_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_src),
    .dev_07_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_priv),
    .dev_07_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_rvso),
    .dev_07_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_07_req_o_fence),
    .dev_08_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_addr),
    .dev_08_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_data),
    .dev_08_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_ben),
    .dev_08_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_stb),
    .dev_08_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_rw),
    .dev_08_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_src),
    .dev_08_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_priv),
    .dev_08_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_rvso),
    .dev_08_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_08_req_o_fence),
    .dev_09_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_addr),
    .dev_09_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_data),
    .dev_09_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_ben),
    .dev_09_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_stb),
    .dev_09_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_rw),
    .dev_09_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_src),
    .dev_09_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_priv),
    .dev_09_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_rvso),
    .dev_09_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_09_req_o_fence),
    .dev_10_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_addr),
    .dev_10_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_data),
    .dev_10_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_ben),
    .dev_10_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_stb),
    .dev_10_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_rw),
    .dev_10_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_src),
    .dev_10_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_priv),
    .dev_10_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_rvso),
    .dev_10_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_10_req_o_fence),
    .dev_11_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_addr),
    .dev_11_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_data),
    .dev_11_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_ben),
    .dev_11_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_stb),
    .dev_11_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_rw),
    .dev_11_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_src),
    .dev_11_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_priv),
    .dev_11_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_rvso),
    .dev_11_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_11_req_o_fence),
    .dev_12_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_addr),
    .dev_12_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_data),
    .dev_12_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_ben),
    .dev_12_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_stb),
    .dev_12_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_rw),
    .dev_12_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_src),
    .dev_12_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_priv),
    .dev_12_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_rvso),
    .dev_12_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_12_req_o_fence),
    .dev_13_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_addr),
    .dev_13_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_data),
    .dev_13_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_ben),
    .dev_13_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_stb),
    .dev_13_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_rw),
    .dev_13_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_src),
    .dev_13_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_priv),
    .dev_13_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_rvso),
    .dev_13_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_13_req_o_fence),
    .dev_14_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_addr),
    .dev_14_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_data),
    .dev_14_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_ben),
    .dev_14_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_stb),
    .dev_14_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_rw),
    .dev_14_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_src),
    .dev_14_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_priv),
    .dev_14_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_rvso),
    .dev_14_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_14_req_o_fence),
    .dev_15_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_addr),
    .dev_15_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_data),
    .dev_15_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_ben),
    .dev_15_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_stb),
    .dev_15_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_rw),
    .dev_15_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_src),
    .dev_15_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_priv),
    .dev_15_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_rvso),
    .dev_15_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_15_req_o_fence),
    .dev_16_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_addr),
    .dev_16_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_data),
    .dev_16_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_ben),
    .dev_16_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_stb),
    .dev_16_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_rw),
    .dev_16_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_src),
    .dev_16_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_priv),
    .dev_16_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_rvso),
    .dev_16_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_16_req_o_fence),
    .dev_17_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_addr),
    .dev_17_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_data),
    .dev_17_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_ben),
    .dev_17_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_stb),
    .dev_17_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_rw),
    .dev_17_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_src),
    .dev_17_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_priv),
    .dev_17_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_rvso),
    .dev_17_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_17_req_o_fence),
    .dev_18_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_addr),
    .dev_18_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_data),
    .dev_18_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_ben),
    .dev_18_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_stb),
    .dev_18_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_rw),
    .dev_18_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_src),
    .dev_18_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_priv),
    .dev_18_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_rvso),
    .dev_18_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_18_req_o_fence),
    .dev_19_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_addr),
    .dev_19_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_data),
    .dev_19_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_ben),
    .dev_19_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_stb),
    .dev_19_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_rw),
    .dev_19_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_src),
    .dev_19_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_priv),
    .dev_19_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_rvso),
    .dev_19_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_19_req_o_fence),
    .dev_20_req_o_addr(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_addr),
    .dev_20_req_o_data(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_data),
    .dev_20_req_o_ben(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_ben),
    .dev_20_req_o_stb(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_stb),
    .dev_20_req_o_rw(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_rw),
    .dev_20_req_o_src(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_src),
    .dev_20_req_o_priv(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_priv),
    .dev_20_req_o_rvso(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_rvso),
    .dev_20_req_o_fence(io_system_neorv32_bus_io_switch_inst_dev_20_req_o_fence));
  assign n477_o = io_req[31:0]; // extract
  assign n478_o = io_req[63:32]; // extract
  assign n479_o = io_req[67:64]; // extract
  assign n480_o = io_req[68]; // extract
  assign n481_o = io_req[69]; // extract
  assign n482_o = io_req[70]; // extract
  assign n483_o = io_req[71]; // extract
  assign n484_o = io_req[72]; // extract
  assign n485_o = io_req[73]; // extract
  assign n486_o = {io_system_neorv32_bus_io_switch_inst_main_rsp_o_err, io_system_neorv32_bus_io_switch_inst_main_rsp_o_ack, io_system_neorv32_bus_io_switch_inst_main_rsp_o_data};
  assign n488_o = {io_system_neorv32_bus_io_switch_inst_dev_00_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_00_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_00_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_00_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_00_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_00_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_00_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_00_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_00_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1056:74  */
  assign n490_o = iodev_rsp[713:680]; // extract
  assign n491_o = n490_o[31:0]; // extract
  assign n492_o = n490_o[32]; // extract
  assign n493_o = n490_o[33]; // extract
  assign n494_o = {io_system_neorv32_bus_io_switch_inst_dev_01_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_01_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_01_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_01_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_01_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_01_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_01_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_01_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_01_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1057:74  */
  assign n496_o = iodev_rsp[679:646]; // extract
  assign n497_o = n496_o[31:0]; // extract
  assign n498_o = n496_o[32]; // extract
  assign n499_o = n496_o[33]; // extract
  assign n500_o = {io_system_neorv32_bus_io_switch_inst_dev_02_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_02_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_02_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_02_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_02_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_02_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_02_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_02_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_02_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1058:74  */
  assign n502_o = iodev_rsp[645:612]; // extract
  assign n503_o = n502_o[31:0]; // extract
  assign n504_o = n502_o[32]; // extract
  assign n505_o = n502_o[33]; // extract
  assign n506_o = {io_system_neorv32_bus_io_switch_inst_dev_03_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_03_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_03_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_03_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_03_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_03_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_03_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_03_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_03_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1059:74  */
  assign n508_o = iodev_rsp[611:578]; // extract
  assign n509_o = n508_o[31:0]; // extract
  assign n510_o = n508_o[32]; // extract
  assign n511_o = n508_o[33]; // extract
  assign n512_o = {io_system_neorv32_bus_io_switch_inst_dev_04_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_04_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_04_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_04_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_04_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_04_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_04_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_04_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_04_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1060:74  */
  assign n514_o = iodev_rsp[577:544]; // extract
  assign n515_o = n514_o[31:0]; // extract
  assign n516_o = n514_o[32]; // extract
  assign n517_o = n514_o[33]; // extract
  assign n518_o = {io_system_neorv32_bus_io_switch_inst_dev_05_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_05_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_05_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_05_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_05_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_05_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_05_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_05_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_05_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1061:74  */
  assign n520_o = iodev_rsp[543:510]; // extract
  assign n521_o = n520_o[31:0]; // extract
  assign n522_o = n520_o[32]; // extract
  assign n523_o = n520_o[33]; // extract
  assign n524_o = {io_system_neorv32_bus_io_switch_inst_dev_06_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_06_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_06_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_06_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_06_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_06_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_06_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_06_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_06_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1062:74  */
  assign n526_o = iodev_rsp[509:476]; // extract
  assign n527_o = n526_o[31:0]; // extract
  assign n528_o = n526_o[32]; // extract
  assign n529_o = n526_o[33]; // extract
  assign n530_o = {io_system_neorv32_bus_io_switch_inst_dev_07_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_07_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_07_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_07_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_07_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_07_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_07_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_07_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_07_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1063:74  */
  assign n532_o = iodev_rsp[475:442]; // extract
  assign n533_o = n532_o[31:0]; // extract
  assign n534_o = n532_o[32]; // extract
  assign n535_o = n532_o[33]; // extract
  assign n536_o = {io_system_neorv32_bus_io_switch_inst_dev_08_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_08_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_08_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_08_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_08_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_08_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_08_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_08_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_08_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1064:74  */
  assign n538_o = iodev_rsp[441:408]; // extract
  assign n539_o = n538_o[31:0]; // extract
  assign n540_o = n538_o[32]; // extract
  assign n541_o = n538_o[33]; // extract
  assign n542_o = {io_system_neorv32_bus_io_switch_inst_dev_09_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_09_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_09_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_09_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_09_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_09_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_09_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_09_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_09_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1065:74  */
  assign n544_o = iodev_rsp[407:374]; // extract
  assign n545_o = n544_o[31:0]; // extract
  assign n546_o = n544_o[32]; // extract
  assign n547_o = n544_o[33]; // extract
  assign n548_o = {io_system_neorv32_bus_io_switch_inst_dev_10_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_10_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_10_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_10_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_10_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_10_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_10_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_10_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_10_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1066:74  */
  assign n550_o = iodev_rsp[373:340]; // extract
  assign n551_o = n550_o[31:0]; // extract
  assign n552_o = n550_o[32]; // extract
  assign n553_o = n550_o[33]; // extract
  assign n554_o = {io_system_neorv32_bus_io_switch_inst_dev_11_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_11_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_11_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_11_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_11_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_11_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_11_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_11_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_11_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1067:74  */
  assign n556_o = iodev_rsp[339:306]; // extract
  assign n557_o = n556_o[31:0]; // extract
  assign n558_o = n556_o[32]; // extract
  assign n559_o = n556_o[33]; // extract
  assign n560_o = {io_system_neorv32_bus_io_switch_inst_dev_12_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_12_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_12_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_12_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_12_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_12_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_12_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_12_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_12_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1068:74  */
  assign n562_o = iodev_rsp[305:272]; // extract
  assign n563_o = n562_o[31:0]; // extract
  assign n564_o = n562_o[32]; // extract
  assign n565_o = n562_o[33]; // extract
  assign n566_o = {io_system_neorv32_bus_io_switch_inst_dev_13_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_13_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_13_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_13_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_13_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_13_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_13_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_13_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_13_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1069:74  */
  assign n568_o = iodev_rsp[271:238]; // extract
  assign n569_o = n568_o[31:0]; // extract
  assign n570_o = n568_o[32]; // extract
  assign n571_o = n568_o[33]; // extract
  assign n572_o = {io_system_neorv32_bus_io_switch_inst_dev_14_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_14_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_14_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_14_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_14_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_14_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_14_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_14_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_14_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1070:74  */
  assign n574_o = iodev_rsp[237:204]; // extract
  assign n575_o = n574_o[31:0]; // extract
  assign n576_o = n574_o[32]; // extract
  assign n577_o = n574_o[33]; // extract
  assign n578_o = {io_system_neorv32_bus_io_switch_inst_dev_15_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_15_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_15_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_15_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_15_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_15_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_15_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_15_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_15_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1071:74  */
  assign n580_o = iodev_rsp[203:170]; // extract
  assign n581_o = n580_o[31:0]; // extract
  assign n582_o = n580_o[32]; // extract
  assign n583_o = n580_o[33]; // extract
  assign n584_o = {io_system_neorv32_bus_io_switch_inst_dev_16_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_16_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_16_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_16_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_16_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_16_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_16_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_16_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_16_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1072:74  */
  assign n586_o = iodev_rsp[169:136]; // extract
  assign n587_o = n586_o[31:0]; // extract
  assign n588_o = n586_o[32]; // extract
  assign n589_o = n586_o[33]; // extract
  assign n590_o = {io_system_neorv32_bus_io_switch_inst_dev_17_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_17_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_17_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_17_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_17_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_17_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_17_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_17_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_17_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1073:74  */
  assign n592_o = iodev_rsp[135:102]; // extract
  assign n593_o = n592_o[31:0]; // extract
  assign n594_o = n592_o[32]; // extract
  assign n595_o = n592_o[33]; // extract
  assign n596_o = {io_system_neorv32_bus_io_switch_inst_dev_18_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_18_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_18_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_18_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_18_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_18_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_18_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_18_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_18_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1074:74  */
  assign n598_o = iodev_rsp[101:68]; // extract
  assign n599_o = n598_o[31:0]; // extract
  assign n600_o = n598_o[32]; // extract
  assign n601_o = n598_o[33]; // extract
  assign n602_o = {io_system_neorv32_bus_io_switch_inst_dev_19_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_19_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_19_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_19_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_19_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_19_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_19_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_19_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_19_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1075:74  */
  assign n604_o = iodev_rsp[67:34]; // extract
  assign n605_o = n604_o[31:0]; // extract
  assign n606_o = n604_o[32]; // extract
  assign n607_o = n604_o[33]; // extract
  assign n608_o = {io_system_neorv32_bus_io_switch_inst_dev_20_req_o_fence, io_system_neorv32_bus_io_switch_inst_dev_20_req_o_rvso, io_system_neorv32_bus_io_switch_inst_dev_20_req_o_priv, io_system_neorv32_bus_io_switch_inst_dev_20_req_o_src, io_system_neorv32_bus_io_switch_inst_dev_20_req_o_rw, io_system_neorv32_bus_io_switch_inst_dev_20_req_o_stb, io_system_neorv32_bus_io_switch_inst_dev_20_req_o_ben, io_system_neorv32_bus_io_switch_inst_dev_20_req_o_data, io_system_neorv32_bus_io_switch_inst_dev_20_req_o_addr};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1076:74  */
  assign n610_o = iodev_rsp[33:0]; // extract
  assign n611_o = n610_o[31:0]; // extract
  assign n612_o = n610_o[32]; // extract
  assign n613_o = n610_o[33]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1199:7  */
  neorv32_mtime io_system_neorv32_mtime_inst_true_neorv32_mtime_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .bus_req_i_addr(n624_o),
    .bus_req_i_data(n625_o),
    .bus_req_i_ben(n626_o),
    .bus_req_i_stb(n627_o),
    .bus_req_i_rw(n628_o),
    .bus_req_i_src(n629_o),
    .bus_req_i_priv(n630_o),
    .bus_req_i_rvso(n631_o),
    .bus_req_i_fence(n632_o),
    .bus_rsp_o_data(io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_data),
    .bus_rsp_o_ack(io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_ack),
    .bus_rsp_o_err(io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_err),
    .time_o(io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_time_o),
    .irq_o(io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_irq_o));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1203:31  */
  assign n623_o = iodev_req[739:666]; // extract
  assign n624_o = n623_o[31:0]; // extract
  assign n625_o = n623_o[63:32]; // extract
  assign n626_o = n623_o[67:64]; // extract
  assign n627_o = n623_o[68]; // extract
  assign n628_o = n623_o[69]; // extract
  assign n629_o = n623_o[70]; // extract
  assign n630_o = n623_o[71]; // extract
  assign n631_o = n623_o[72]; // extract
  assign n632_o = n623_o[73]; // extract
  assign n633_o = {io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_err, io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_ack, io_system_neorv32_mtime_inst_true_neorv32_mtime_inst_bus_rsp_o_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1212:22  */
  assign n638_o = ~rstn_sys;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1215:50  */
  assign n641_o = mtime_time[31:0]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1220:47  */
  assign n646_o = mtime_time[63:32]; // extract
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1587:5  */
  neorv32_sysinfo_0_16384_8192_4_4_64_4_64_32_32_8_256_ad514a383a71baac85f4c0ffc48c0bd10a15d22b io_system_neorv32_sysinfo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .bus_req_i_addr(n684_o),
    .bus_req_i_data(n685_o),
    .bus_req_i_ben(n686_o),
    .bus_req_i_stb(n687_o),
    .bus_req_i_rw(n688_o),
    .bus_req_i_src(n689_o),
    .bus_req_i_priv(n690_o),
    .bus_req_i_rvso(n691_o),
    .bus_req_i_fence(n692_o),
    .bus_rsp_o_data(io_system_neorv32_sysinfo_inst_bus_rsp_o_data),
    .bus_rsp_o_ack(io_system_neorv32_sysinfo_inst_bus_rsp_o_ack),
    .bus_rsp_o_err(io_system_neorv32_sysinfo_inst_bus_rsp_o_err));
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1634:29  */
  assign n683_o = iodev_req[1479:1406]; // extract
  assign n684_o = n683_o[31:0]; // extract
  assign n685_o = n683_o[63:32]; // extract
  assign n686_o = n683_o[67:64]; // extract
  assign n687_o = n683_o[68]; // extract
  assign n688_o = n683_o[69]; // extract
  assign n689_o = n683_o[70]; // extract
  assign n690_o = n683_o[71]; // extract
  assign n691_o = n683_o[72]; // extract
  assign n692_o = n683_o[73]; // extract
  assign n693_o = {io_system_neorv32_sysinfo_inst_bus_rsp_o_err, io_system_neorv32_sysinfo_inst_bus_rsp_o_ack, io_system_neorv32_sysinfo_inst_bus_rsp_o_data};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:430:7  */
  always @(negedge clk_i or posedge n197_o)
    if (n197_o)
      n697_q <= 4'b0000;
    else
      n697_q <= n225_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:430:7  */
  always @(negedge clk_i or posedge n197_o)
    if (n197_o)
      n699_q <= 1'b0;
    else
      n699_q <= n241_o;
  assign n713_o = {n488_o, n494_o, n500_o, n506_o, n512_o, n518_o, n524_o, n530_o, n536_o, n542_o, n548_o, n554_o, n560_o, n566_o, n572_o, n578_o, n584_o, n590_o, n596_o, n602_o, n608_o};
  assign n714_o = {34'b0000000000000000000000000000000000, n693_o, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, n633_o, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000};
  assign n715_o = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  assign n716_o = {n365_o, n364_o, n363_o, n362_o, n361_o, n360_o, n359_o, n358_o, n357_o, n356_o, n355_o, n354_o, n353_o, n352_o, n351_o, n350_o};
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1214:9  */
  always @(posedge clk_i or posedge n638_o)
    if (n638_o)
      n717_q <= 32'b00000000000000000000000000000000;
    else
      n717_q <= n641_o;
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_top.vhd:1212:9  */
  assign n718_o = {n646_o, n717_q};
endmodule

module neorv32_litex_core_complex
  (input  clk_i,
   input  rstn_i,
   input  jtag_trst_i,
   input  jtag_tck_i,
   input  jtag_tdi_i,
   input  jtag_tms_i,
   input  [31:0] wb_dat_i,
   input  wb_ack_i,
   input  wb_err_i,
   input  mext_irq_i,
   output jtag_tdo_o,
   output [31:0] wb_adr_o,
   output [31:0] wb_dat_o,
   output wb_we_o,
   output [3:0] wb_sel_o,
   output wb_stb_o,
   output wb_cyc_o);
  wire neorv32_core_complex_n7;
  wire [31:0] neorv32_core_complex_n8;
  wire [31:0] neorv32_core_complex_n9;
  wire neorv32_core_complex_n10;
  wire [3:0] neorv32_core_complex_n11;
  wire neorv32_core_complex_n12;
  wire neorv32_core_complex_n13;
  localparam [31:0] n14_o = 32'b00000000000000000000000000000000;
  localparam n15_o = 1'b0;
  localparam n16_o = 1'b0;
  localparam n21_o = 1'b0;
  localparam n24_o = 1'b0;
  localparam [63:0] n27_o = 64'b0000000000000000000000000000000000000000000000000000000000000000;
  localparam n29_o = 1'b0;
  localparam n31_o = 1'b0;
  localparam n33_o = 1'b0;
  localparam n35_o = 1'b0;
  localparam n38_o = 1'b0;
  localparam n40_o = 1'b0;
  localparam n42_o = 1'b0;
  localparam n43_o = 1'b1;
  localparam n44_o = 1'b1;
  localparam n46_o = 1'b1;
  localparam n48_o = 1'b1;
  localparam [31:0] n51_o = 32'b00000000000000000000000000000000;
  localparam n55_o = 1'b0;
  localparam [31:0] n56_o = 32'b00000000000000000000000000000000;
  localparam n57_o = 1'b0;
  localparam n58_o = 1'b0;
  wire neorv32_core_complex_jtag_tdo_o;
  wire [31:0] neorv32_core_complex_xbus_adr_o;
  wire [31:0] neorv32_core_complex_xbus_dat_o;
  wire neorv32_core_complex_xbus_we_o;
  wire [3:0] neorv32_core_complex_xbus_sel_o;
  wire neorv32_core_complex_xbus_stb_o;
  wire neorv32_core_complex_xbus_cyc_o;
  wire neorv32_core_complex_slink_rx_rdy_o;
  wire [31:0] neorv32_core_complex_slink_tx_dat_o;
  wire neorv32_core_complex_slink_tx_val_o;
  wire neorv32_core_complex_slink_tx_lst_o;
  wire neorv32_core_complex_xip_csn_o;
  wire neorv32_core_complex_xip_clk_o;
  wire neorv32_core_complex_xip_dat_o;
  wire [63:0] neorv32_core_complex_gpio_o;
  wire neorv32_core_complex_uart0_txd_o;
  wire neorv32_core_complex_uart0_rts_o;
  wire neorv32_core_complex_uart1_txd_o;
  wire neorv32_core_complex_uart1_rts_o;
  wire neorv32_core_complex_spi_clk_o;
  wire neorv32_core_complex_spi_dat_o;
  wire [7:0] neorv32_core_complex_spi_csn_o;
  wire neorv32_core_complex_sdi_dat_o;
  wire neorv32_core_complex_twi_sda_o;
  wire neorv32_core_complex_twi_scl_o;
  wire neorv32_core_complex_onewire_o;
  wire [11:0] neorv32_core_complex_pwm_o;
  wire [31:0] neorv32_core_complex_cfs_out_o;
  wire neorv32_core_complex_neoled_o;
  wire [63:0] neorv32_core_complex_mtime_time_o;
  assign jtag_tdo_o = neorv32_core_complex_n7; //(module output)
  assign wb_adr_o = neorv32_core_complex_n8; //(module output)
  assign wb_dat_o = neorv32_core_complex_n9; //(module output)
  assign wb_we_o = neorv32_core_complex_n10; //(module output)
  assign wb_sel_o = neorv32_core_complex_n11; //(module output)
  assign wb_stb_o = neorv32_core_complex_n12; //(module output)
  assign wb_cyc_o = neorv32_core_complex_n13; //(module output)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_litex_core_complex.vhd:201:20  */
  assign neorv32_core_complex_n7 = neorv32_core_complex_jtag_tdo_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_litex_core_complex.vhd:204:20  */
  assign neorv32_core_complex_n8 = neorv32_core_complex_xbus_adr_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_litex_core_complex.vhd:206:20  */
  assign neorv32_core_complex_n9 = neorv32_core_complex_xbus_dat_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_litex_core_complex.vhd:207:20  */
  assign neorv32_core_complex_n10 = neorv32_core_complex_xbus_we_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_litex_core_complex.vhd:208:20  */
  assign neorv32_core_complex_n11 = neorv32_core_complex_xbus_sel_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_litex_core_complex.vhd:209:20  */
  assign neorv32_core_complex_n12 = neorv32_core_complex_xbus_stb_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_litex_core_complex.vhd:210:20  */
  assign neorv32_core_complex_n13 = neorv32_core_complex_xbus_cyc_o; // (signal)
  /* /home/micko/src/litex/litex/litex/soc/cores/cpu/neorv32/neorv32_litex_core_complex.vhd:158:3  */
  neorv32_top_0_0_4_0_64_4_16384_8192_4_64_4_64_1024_32_32_8_256_0_0_1_1_1_1_1_1_0_1_32_32_1_1_1_ba529af7aa7a6f941b636046ab20a941c3aa1b01 neorv32_core_complex (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .jtag_trst_i(jtag_trst_i),
    .jtag_tck_i(jtag_tck_i),
    .jtag_tdi_i(jtag_tdi_i),
    .jtag_tms_i(jtag_tms_i),
    .xbus_dat_i(wb_dat_i),
    .xbus_ack_i(wb_ack_i),
    .xbus_err_i(wb_err_i),
    .slink_rx_dat_i(n14_o),
    .slink_rx_val_i(n15_o),
    .slink_rx_lst_i(n16_o),
    .slink_tx_rdy_i(n21_o),
    .xip_dat_i(n24_o),
    .gpio_i(n27_o),
    .uart0_rxd_i(n29_o),
    .uart0_cts_i(n31_o),
    .uart1_rxd_i(n33_o),
    .uart1_cts_i(n35_o),
    .spi_dat_i(n38_o),
    .sdi_clk_i(n40_o),
    .sdi_dat_i(n42_o),
    .sdi_csn_i(n43_o),
    .twi_sda_i(n44_o),
    .twi_scl_i(n46_o),
    .onewire_i(n48_o),
    .cfs_in_i(n51_o),
    .gptmr_trig_i(n55_o),
    .xirq_i(n56_o),
    .mtime_irq_i(n57_o),
    .msw_irq_i(n58_o),
    .mext_irq_i(mext_irq_i),
    .jtag_tdo_o(neorv32_core_complex_jtag_tdo_o),
    .xbus_adr_o(neorv32_core_complex_xbus_adr_o),
    .xbus_dat_o(neorv32_core_complex_xbus_dat_o),
    .xbus_we_o(neorv32_core_complex_xbus_we_o),
    .xbus_sel_o(neorv32_core_complex_xbus_sel_o),
    .xbus_stb_o(neorv32_core_complex_xbus_stb_o),
    .xbus_cyc_o(neorv32_core_complex_xbus_cyc_o),
    .slink_rx_rdy_o(),
    .slink_tx_dat_o(),
    .slink_tx_val_o(),
    .slink_tx_lst_o(),
    .xip_csn_o(),
    .xip_clk_o(),
    .xip_dat_o(),
    .gpio_o(),
    .uart0_txd_o(),
    .uart0_rts_o(),
    .uart1_txd_o(),
    .uart1_rts_o(),
    .spi_clk_o(),
    .spi_dat_o(),
    .spi_csn_o(),
    .sdi_dat_o(),
    .twi_sda_o(),
    .twi_scl_o(),
    .onewire_o(),
    .pwm_o(),
    .cfs_out_o(),
    .neoled_o(),
    .mtime_time_o());
endmodule

